// key=00

module s27_obf(CK, G0, G1, G2, G3, G17, keyinput);
input CK;
input G0;
input G1;
input G2;
input G3;
input [1:0] keyinput;
output G17;
wire G5;
wire G6;
wire G7;
wire G14;
wire G8;
wire G15;
wire G16;
wire G9;
wire G10;
wire G12;
wire G13;
wire G13_obf;
wire G11;
wire G11_obf;
dff DFF_0(CK, G5, G10);
dff DFF_1(CK, G6, G11);
dff DFF_2(CK, G7, G13);
not NOT_0(G14, G0);
not NOT_1(G17, G11);
and AND2_0(G8, G14, G6);
or OR2_0(G15, G12, G8);
or OR2_1(G16, G3, G8);
nand NAND2_0(G9, G16, G15);
nor NOR2_0(G10, G14, G11);
nor NOR2_2(G12, G1, G7);
xor tag0(G13, keyinput[0], G13_obf);
nor NOR2_3(G13_obf, G2, G12);
xor tag1(G11, keyinput[1], G11_obf);
nor NOR2_1(G11_obf, G5, G9);
endmodule