module c6288(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,
  G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G4,G5,G6,G6257,G6258,G6259,G6260,
  G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,
  G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,G6281,G6282,G6283,G6284,
  G6285,G6286,G6287,G6288,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32;
output G6257,G6258,G6259,G6260,G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,
  G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
  G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288;

  wire G545,G548,G551,G554,G557,G560,G563,G566,G569,G572,G575,G578,G581,G584,
    G587,G590,G593,G596,G599,G602,G605,G608,G611,G614,G617,G620,G623,G626,G629,
    G632,G635,G638,G641,G644,G647,G650,G653,G656,G659,G662,G665,G668,G671,G674,
    G677,G680,G683,G686,G689,G692,G695,G698,G701,G704,G707,G710,G713,G716,G719,
    G722,G725,G728,G731,G734,G737,G740,G743,G746,G749,G752,G755,G758,G761,G764,
    G767,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,G809,
    G812,G815,G818,G821,G824,G827,G830,G833,G836,G839,G842,G845,G848,G851,G854,
    G857,G860,G863,G866,G869,G872,G875,G878,G881,G884,G887,G890,G893,G896,G899,
    G902,G905,G908,G911,G914,G917,G920,G923,G926,G929,G932,G935,G938,G941,G944,
    G947,G950,G953,G956,G959,G962,G965,G968,G971,G974,G977,G980,G983,G986,G989,
    G992,G995,G998,G1001,G1004,G1007,G1010,G1013,G1016,G1019,G1022,G1025,G1028,
    G1031,G1034,G1037,G1040,G1043,G1046,G1049,G1052,G1055,G1058,G1061,G1064,
    G1067,G1070,G1073,G1076,G1079,G1082,G1085,G1088,G1091,G1094,G1097,G1100,
    G1103,G1106,G1109,G1112,G1115,G1118,G1121,G1124,G1127,G1130,G1133,G1136,
    G1139,G1142,G1145,G1148,G1151,G1154,G1157,G1160,G1163,G1166,G1169,G1172,
    G1175,G1178,G1181,G1184,G1187,G1190,G1193,G1196,G1199,G1202,G1205,G1208,
    G1211,G1214,G1217,G1220,G1223,G1226,G1229,G1232,G1235,G1238,G1241,G1244,
    G1247,G1250,G1253,G1256,G1259,G1262,G1265,G1268,G1271,G1274,G1277,G1280,
    G1283,G1286,G1289,G1292,G1295,G1298,G1301,G1304,G1307,G1310,G1314,G1318,
    G1322,G1326,G1330,G1334,G1338,G1342,G1346,G1350,G1354,G1358,G1362,G1366,
    G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,G1381,
    G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,
    G1394,G1395,G1396,G1397,G1398,G1399,G1400,G1403,G1406,G1409,G1412,G1415,
    G1418,G1421,G1424,G1427,G1430,G1433,G1436,G1439,G1442,G1445,G1449,G1453,
    G1457,G1461,G1465,G1469,G1473,G1477,G1481,G1485,G1489,G1493,G1497,G1501,
    G1505,G1506,G1507,G1510,G1511,G1512,G1515,G1516,G1517,G1520,G1521,G1522,
    G1525,G1526,G1527,G1530,G1531,G1532,G1535,G1536,G1537,G1540,G1541,G1542,
    G1545,G1546,G1547,G1550,G1551,G1552,G1555,G1556,G1557,G1560,G1561,G1562,
    G1565,G1566,G1567,G1570,G1571,G1572,G1575,G1576,G1577,G1580,G1583,G1586,
    G1589,G1592,G1595,G1598,G1601,G1604,G1607,G1610,G1613,G1616,G1619,G1622,
    G1626,G1630,G1634,G1638,G1642,G1646,G1650,G1654,G1658,G1662,G1666,G1670,
    G1674,G1678,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,
    G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,G1701,G1702,G1703,
    G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1715,G1718,G1721,
    G1724,G1727,G1730,G1733,G1736,G1739,G1742,G1745,G1748,G1751,G1754,G1757,
    G1761,G1765,G1769,G1773,G1777,G1781,G1785,G1789,G1793,G1797,G1801,G1805,
    G1809,G1813,G1817,G1818,G1819,G1822,G1823,G1824,G1827,G1828,G1829,G1832,
    G1833,G1834,G1837,G1838,G1839,G1842,G1843,G1844,G1847,G1848,G1849,G1852,
    G1853,G1854,G1857,G1858,G1859,G1862,G1863,G1864,G1867,G1868,G1869,G1872,
    G1873,G1874,G1877,G1878,G1879,G1882,G1883,G1884,G1887,G1888,G1889,G1892,
    G1895,G1899,G1902,G1905,G1908,G1911,G1914,G1917,G1920,G1923,G1926,G1929,
    G1932,G1935,G1938,G1942,G1943,G1944,G1948,G1952,G1956,G1960,G1964,G1968,
    G1972,G1976,G1980,G1984,G1988,G1992,G1996,G1997,G1998,G2001,G2002,G2003,
    G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,
    G2016,G2017,G2018,G2019,G2020,G2021,G2022,G2023,G2024,G2025,G2026,G2027,
    G2030,G2034,G2037,G2040,G2043,G2046,G2049,G2052,G2055,G2058,G2061,G2064,
    G2067,G2070,G2073,G2077,G2078,G2079,G2082,G2086,G2090,G2094,G2098,G2102,
    G2106,G2110,G2114,G2118,G2122,G2126,G2130,G2134,G2135,G2136,G2139,G2142,
    G2146,G2147,G2148,G2151,G2152,G2153,G2156,G2157,G2158,G2161,G2162,G2163,
    G2166,G2167,G2168,G2171,G2172,G2173,G2176,G2177,G2178,G2181,G2182,G2183,
    G2186,G2187,G2188,G2191,G2192,G2193,G2196,G2197,G2198,G2201,G2202,G2203,
    G2206,G2207,G2208,G2211,G2214,G2218,G2219,G2220,G2223,G2226,G2229,G2232,
    G2235,G2238,G2241,G2244,G2247,G2250,G2253,G2256,G2260,G2261,G2262,G2265,
    G2269,G2273,G2277,G2281,G2285,G2289,G2293,G2297,G2301,G2305,G2309,G2313,
    G2314,G2315,G2318,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,
    G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,G2341,G2342,
    G2343,G2344,G2345,G2346,G2349,G2353,G2354,G2355,G2358,G2361,G2364,G2367,
    G2370,G2373,G2376,G2379,G2382,G2385,G2388,G2391,G2394,G2398,G2399,G2400,
    G2403,G2406,G2410,G2414,G2418,G2422,G2426,G2430,G2434,G2438,G2442,G2446,
    G2450,G2454,G2458,G2459,G2460,G2463,G2466,G2470,G2471,G2472,G2473,G2474,
    G2477,G2478,G2479,G2482,G2483,G2484,G2487,G2488,G2489,G2492,G2493,G2494,
    G2497,G2498,G2499,G2502,G2503,G2504,G2507,G2508,G2509,G2512,G2513,G2514,
    G2517,G2518,G2519,G2522,G2523,G2524,G2527,G2528,G2529,G2532,G2535,G2539,
    G2540,G2541,G2544,G2547,G2550,G2553,G2556,G2559,G2562,G2565,G2568,G2571,
    G2574,G2577,G2581,G2582,G2583,G2586,G2590,G2594,G2598,G2602,G2606,G2610,
    G2614,G2618,G2622,G2626,G2630,G2634,G2635,G2636,G2639,G2643,G2644,G2645,
    G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,
    G2660,G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2673,
    G2677,G2678,G2679,G2682,G2685,G2689,G2692,G2695,G2698,G2701,G2704,G2707,
    G2710,G2713,G2716,G2719,G2722,G2726,G2727,G2728,G2731,G2734,G2738,G2739,
    G2740,G2744,G2748,G2752,G2756,G2760,G2764,G2768,G2772,G2776,G2780,G2784,
    G2785,G2786,G2789,G2792,G2796,G2797,G2798,G2801,G2802,G2803,G2806,G2807,
    G2808,G2811,G2812,G2813,G2816,G2817,G2818,G2821,G2822,G2823,G2826,G2827,
    G2828,G2831,G2832,G2833,G2836,G2837,G2838,G2841,G2842,G2843,G2846,G2847,
    G2848,G2851,G2852,G2853,G2856,G2859,G2863,G2864,G2865,G2868,G2872,G2875,
    G2878,G2881,G2884,G2887,G2890,G2893,G2896,G2899,G2902,G2906,G2907,G2908,
    G2911,G2915,G2916,G2917,G2920,G2924,G2928,G2932,G2936,G2940,G2944,G2948,
    G2952,G2956,G2960,G2961,G2962,G2965,G2969,G2970,G2971,G2974,G2977,G2981,
    G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,
    G2994,G2995,G2996,G2997,G2998,G2999,G3000,G3001,G3004,G3008,G3009,G3010,
    G3013,G3016,G3020,G3021,G3022,G3025,G3028,G3031,G3034,G3037,G3040,G3043,
    G3046,G3049,G3052,G3056,G3057,G3058,G3061,G3064,G3068,G3069,G3070,G3073,
    G3077,G3081,G3085,G3089,G3093,G3097,G3101,G3105,G3109,G3113,G3114,G3115,
    G3118,G3121,G3125,G3126,G3127,G3130,G3134,G3135,G3136,G3139,G3140,G3141,
    G3144,G3145,G3146,G3149,G3150,G3151,G3154,G3155,G3156,G3159,G3160,G3161,
    G3164,G3165,G3166,G3169,G3170,G3171,G3174,G3175,G3176,G3179,G3180,G3181,
    G3184,G3187,G3191,G3192,G3193,G3196,G3200,G3201,G3202,G3205,G3208,G3211,
    G3214,G3217,G3220,G3223,G3226,G3229,G3232,G3236,G3237,G3238,G3241,G3245,
    G3246,G3247,G3250,G3253,G3257,G3261,G3265,G3269,G3273,G3277,G3281,G3285,
    G3289,G3293,G3294,G3295,G3298,G3302,G3303,G3304,G3307,G3310,G3314,G3315,
    G3316,G3317,G3318,G3319,G3320,G3321,G3322,G3323,G3324,G3325,G3326,G3327,
    G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3337,G3341,G3342,G3343,G3346,
    G3349,G3353,G3354,G3355,G3358,G3361,G3364,G3367,G3370,G3373,G3376,G3379,
    G3382,G3385,G3389,G3390,G3391,G3394,G3397,G3401,G3402,G3403,G3406,G3410,
    G3414,G3418,G3422,G3426,G3430,G3434,G3438,G3442,G3446,G3447,G3448,G3451,
    G3454,G3458,G3459,G3460,G3463,G3467,G3468,G3469,G3472,G3473,G3474,G3477,
    G3478,G3479,G3482,G3483,G3484,G3487,G3488,G3489,G3492,G3493,G3494,G3497,
    G3498,G3499,G3502,G3503,G3504,G3507,G3508,G3509,G3512,G3513,G3514,G3517,
    G3520,G3524,G3525,G3526,G3529,G3533,G3534,G3535,G3538,G3541,G3545,G3548,
    G3551,G3554,G3557,G3560,G3563,G3566,G3569,G3573,G3574,G3575,G3578,G3582,
    G3583,G3584,G3587,G3590,G3594,G3595,G3596,G3600,G3604,G3608,G3612,G3616,
    G3620,G3624,G3628,G3629,G3630,G3633,G3637,G3638,G3639,G3642,G3645,G3649,
    G3650,G3651,G3654,G3655,G3656,G3657,G3658,G3659,G3660,G3661,G3662,G3663,
    G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3673,G3677,G3678,G3679,G3682,
    G3685,G3689,G3690,G3691,G3694,G3698,G3701,G3704,G3707,G3710,G3713,G3716,
    G3719,G3722,G3726,G3727,G3728,G3731,G3734,G3738,G3739,G3740,G3743,G3747,
    G3748,G3749,G3752,G3756,G3760,G3764,G3768,G3772,G3776,G3780,G3784,G3785,
    G3786,G3789,G3792,G3796,G3797,G3798,G3801,G3805,G3806,G3807,G3810,G3813,
    G3817,G3818,G3819,G3822,G3823,G3824,G3827,G3828,G3829,G3832,G3833,G3834,
    G3837,G3838,G3839,G3842,G3843,G3844,G3847,G3848,G3849,G3852,G3853,G3854,
    G3857,G3860,G3864,G3865,G3866,G3869,G3873,G3874,G3875,G3878,G3881,G3885,
    G3886,G3887,G3890,G3893,G3896,G3899,G3902,G3905,G3908,G3912,G3913,G3914,
    G3917,G3921,G3922,G3923,G3926,G3929,G3933,G3934,G3935,G3938,G3942,G3946,
    G3950,G3954,G3958,G3962,G3966,G3967,G3968,G3971,G3975,G3976,G3977,G3980,
    G3983,G3987,G3988,G3989,G3992,G3996,G3997,G3998,G3999,G4000,G4001,G4002,
    G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4013,G4017,G4018,G4019,
    G4022,G4025,G4029,G4030,G4031,G4034,G4038,G4039,G4040,G4043,G4046,G4049,
    G4052,G4055,G4058,G4061,G4064,G4068,G4069,G4070,G4073,G4076,G4080,G4081,
    G4082,G4085,G4089,G4090,G4091,G4094,G4097,G4101,G4105,G4109,G4113,G4117,
    G4121,G4125,G4129,G4130,G4131,G4134,G4137,G4141,G4142,G4143,G4146,G4150,
    G4151,G4152,G4155,G4158,G4162,G4163,G4164,G4165,G4166,G4169,G4170,G4171,
    G4174,G4175,G4176,G4179,G4180,G4181,G4184,G4185,G4186,G4189,G4190,G4191,
    G4194,G4195,G4196,G4199,G4202,G4206,G4207,G4208,G4211,G4215,G4216,G4217,
    G4220,G4223,G4227,G4228,G4229,G4232,G4235,G4238,G4241,G4244,G4247,G4250,
    G4254,G4255,G4256,G4259,G4263,G4264,G4265,G4268,G4271,G4275,G4276,G4277,
    G4280,G4284,G4288,G4292,G4296,G4300,G4304,G4308,G4309,G4310,G4313,G4317,
    G4318,G4319,G4322,G4325,G4329,G4330,G4331,G4334,G4338,G4339,G4340,G4343,
    G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,
    G4358,G4362,G4363,G4364,G4367,G4370,G4374,G4375,G4376,G4379,G4383,G4384,
    G4385,G4388,G4391,G4395,G4398,G4401,G4404,G4407,G4410,G4413,G4417,G4418,
    G4419,G4422,G4425,G4429,G4430,G4431,G4434,G4438,G4439,G4440,G4443,G4446,
    G4450,G4451,G4452,G4456,G4460,G4464,G4468,G4472,G4476,G4477,G4478,G4481,
    G4484,G4488,G4489,G4490,G4493,G4497,G4498,G4499,G4502,G4505,G4509,G4510,
    G4511,G4514,G4515,G4516,G4519,G4520,G4521,G4524,G4525,G4526,G4529,G4530,
    G4531,G4534,G4535,G4536,G4539,G4540,G4541,G4544,G4547,G4551,G4552,G4553,
    G4556,G4560,G4561,G4562,G4565,G4568,G4572,G4573,G4574,G4577,G4581,G4584,
    G4587,G4590,G4593,G4596,G4600,G4601,G4602,G4605,G4609,G4610,G4611,G4614,
    G4617,G4621,G4622,G4623,G4626,G4630,G4631,G4632,G4635,G4639,G4643,G4647,
    G4651,G4655,G4656,G4657,G4660,G4664,G4665,G4666,G4669,G4672,G4676,G4677,
    G4678,G4681,G4685,G4686,G4687,G4690,G4693,G4697,G4698,G4699,G4700,G4701,
    G4702,G4703,G4704,G4705,G4706,G4707,G4710,G4714,G4715,G4716,G4719,G4722,
    G4726,G4727,G4728,G4731,G4735,G4736,G4737,G4740,G4743,G4747,G4748,G4749,
    G4752,G4755,G4758,G4761,G4764,G4768,G4769,G4770,G4773,G4776,G4780,G4781,
    G4782,G4785,G4789,G4790,G4791,G4794,G4797,G4801,G4802,G4803,G4806,G4810,
    G4814,G4818,G4822,G4826,G4827,G4828,G4831,G4834,G4838,G4839,G4840,G4843,
    G4847,G4848,G4849,G4852,G4855,G4859,G4860,G4861,G4864,G4868,G4869,G4870,
    G4873,G4874,G4875,G4878,G4879,G4880,G4883,G4884,G4885,G4888,G4889,G4890,
    G4893,G4896,G4900,G4901,G4902,G4905,G4909,G4910,G4911,G4914,G4917,G4921,
    G4922,G4923,G4926,G4930,G4931,G4932,G4935,G4938,G4941,G4944,G4947,G4951,
    G4952,G4953,G4956,G4960,G4961,G4962,G4965,G4968,G4972,G4973,G4974,G4977,
    G4981,G4982,G4983,G4986,G4989,G4993,G4997,G5001,G5005,G5009,G5010,G5011,
    G5014,G5018,G5019,G5020,G5023,G5026,G5030,G5031,G5032,G5035,G5039,G5040,
    G5041,G5044,G5047,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,
    G5060,G5061,G5064,G5068,G5069,G5070,G5073,G5076,G5080,G5081,G5082,G5085,
    G5089,G5090,G5091,G5094,G5097,G5101,G5102,G5103,G5106,G5109,G5112,G5115,
    G5118,G5122,G5123,G5124,G5127,G5130,G5134,G5135,G5136,G5139,G5143,G5144,
    G5145,G5148,G5151,G5155,G5156,G5157,G5160,G5164,G5168,G5172,G5176,G5180,
    G5181,G5182,G5185,G5188,G5192,G5193,G5194,G5197,G5201,G5202,G5203,G5206,
    G5209,G5213,G5214,G5215,G5218,G5222,G5223,G5224,G5227,G5228,G5229,G5232,
    G5233,G5234,G5237,G5238,G5239,G5242,G5243,G5244,G5247,G5250,G5254,G5255,
    G5256,G5259,G5263,G5264,G5265,G5268,G5271,G5275,G5276,G5277,G5280,G5284,
    G5285,G5286,G5289,G5292,G5296,G5299,G5302,G5305,G5309,G5310,G5311,G5314,
    G5318,G5319,G5320,G5323,G5326,G5330,G5331,G5332,G5335,G5339,G5340,G5341,
    G5344,G5347,G5351,G5352,G5353,G5357,G5361,G5365,G5366,G5367,G5370,G5374,
    G5375,G5376,G5379,G5382,G5386,G5387,G5388,G5391,G5395,G5396,G5397,G5400,
    G5403,G5407,G5408,G5409,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5421,
    G5425,G5426,G5427,G5430,G5433,G5437,G5438,G5439,G5442,G5446,G5447,G5448,
    G5451,G5454,G5458,G5459,G5460,G5463,G5467,G5470,G5473,G5476,G5480,G5481,
    G5482,G5485,G5488,G5492,G5493,G5494,G5497,G5501,G5502,G5503,G5506,G5509,
    G5513,G5514,G5515,G5518,G5522,G5523,G5524,G5527,G5531,G5535,G5539,G5540,
    G5541,G5544,G5547,G5551,G5552,G5553,G5556,G5560,G5561,G5562,G5565,G5568,
    G5572,G5573,G5574,G5577,G5581,G5582,G5583,G5586,G5589,G5593,G5594,G5595,
    G5598,G5599,G5600,G5603,G5604,G5605,G5608,G5611,G5615,G5616,G5617,G5620,
    G5624,G5625,G5626,G5629,G5632,G5636,G5637,G5638,G5641,G5645,G5646,G5647,
    G5650,G5653,G5657,G5658,G5659,G5662,G5665,G5669,G5670,G5671,G5674,G5678,
    G5679,G5680,G5683,G5686,G5690,G5691,G5692,G5695,G5699,G5700,G5701,G5704,
    G5707,G5711,G5712,G5713,G5716,G5720,G5724,G5725,G5726,G5729,G5733,G5734,
    G5735,G5738,G5741,G5745,G5746,G5747,G5750,G5754,G5755,G5756,G5759,G5762,
    G5766,G5767,G5768,G5771,G5772,G5773,G5774,G5775,G5778,G5782,G5783,G5784,
    G5787,G5790,G5794,G5795,G5796,G5799,G5803,G5804,G5805,G5808,G5811,G5815,
    G5816,G5817,G5820,G5823,G5826,G5830,G5831,G5832,G5835,G5838,G5842,G5843,
    G5844,G5847,G5851,G5852,G5853,G5856,G5859,G5863,G5864,G5865,G5868,G5872,
    G5876,G5877,G5878,G5881,G5884,G5888,G5889,G5890,G5893,G5897,G5898,G5899,
    G5902,G5905,G5909,G5910,G5911,G5914,G5915,G5916,G5919,G5920,G5921,G5924,
    G5927,G5931,G5932,G5933,G5936,G5940,G5941,G5942,G5945,G5948,G5952,G5953,
    G5954,G5957,G5960,G5964,G5965,G5966,G5969,G5973,G5974,G5975,G5978,G5981,
    G5985,G5986,G5987,G5990,G5994,G5995,G5996,G5999,G6003,G6004,G6005,G6008,
    G6011,G6015,G6016,G6017,G6020,G6021,G6022,G6025,G6029,G6030,G6031,G6034,
    G6037,G6041,G6042,G6043,G6046,G6049,G6053,G6054,G6055,G6058,G6061,G6065,
    G6066,G6067,G6070,G6074,G6075,G6076,G6079,G6082,G6086,G6087,G6088,G6091,
    G6092,G6093,G6096,G6099,G6103,G6104,G6105,G6108,G6112,G6113,G6114,G6117,
    G6118,G6119,G6122,G6125,G6129,G6130,G6131,G6134,G6138,G6139,G6140,G6143,
    G6147,G6148,G6149,G6152,G6156,G6157,G6158,G6161,G6165,G6166,G6167,G6170,
    G6174,G6175,G6176,G6179,G6183,G6184,G6185,G6188,G6192,G6193,G6194,G6197,
    G6201,G6202,G6203,G6206,G6210,G6211,G6212,G6215,G6219,G6220,G6221,G6224,
    G6228,G6229,G6230,G6233,G6237,G6238,G6239,G6242,G6246,G6247,G6248,G6251,
    G6255,G6256;

  and AND2_0(G545,G1,G18);
  and AND2_1(G548,G1,G19);
  and AND2_2(G551,G1,G20);
  and AND2_3(G554,G1,G21);
  and AND2_4(G557,G1,G22);
  and AND2_5(G560,G1,G23);
  and AND2_6(G563,G1,G24);
  and AND2_7(G566,G1,G25);
  and AND2_8(G569,G1,G26);
  and AND2_9(G572,G1,G27);
  and AND2_10(G575,G1,G28);
  and AND2_11(G578,G1,G29);
  and AND2_12(G581,G1,G30);
  and AND2_13(G584,G1,G31);
  and AND2_14(G587,G1,G32);
  and AND2_15(G590,G2,G17);
  and AND2_16(G593,G2,G18);
  and AND2_17(G596,G2,G19);
  and AND2_18(G599,G2,G20);
  and AND2_19(G602,G2,G21);
  and AND2_20(G605,G2,G22);
  and AND2_21(G608,G2,G23);
  and AND2_22(G611,G2,G24);
  and AND2_23(G614,G2,G25);
  and AND2_24(G617,G2,G26);
  and AND2_25(G620,G2,G27);
  and AND2_26(G623,G2,G28);
  and AND2_27(G626,G2,G29);
  and AND2_28(G629,G2,G30);
  and AND2_29(G632,G2,G31);
  and AND2_30(G635,G2,G32);
  and AND2_31(G638,G3,G17);
  and AND2_32(G641,G3,G18);
  and AND2_33(G644,G3,G19);
  and AND2_34(G647,G3,G20);
  and AND2_35(G650,G3,G21);
  and AND2_36(G653,G3,G22);
  and AND2_37(G656,G3,G23);
  and AND2_38(G659,G3,G24);
  and AND2_39(G662,G3,G25);
  and AND2_40(G665,G3,G26);
  and AND2_41(G668,G3,G27);
  and AND2_42(G671,G3,G28);
  and AND2_43(G674,G3,G29);
  and AND2_44(G677,G3,G30);
  and AND2_45(G680,G3,G31);
  and AND2_46(G683,G3,G32);
  and AND2_47(G686,G4,G17);
  and AND2_48(G689,G4,G18);
  and AND2_49(G692,G4,G19);
  and AND2_50(G695,G4,G20);
  and AND2_51(G698,G4,G21);
  and AND2_52(G701,G4,G22);
  and AND2_53(G704,G4,G23);
  and AND2_54(G707,G4,G24);
  and AND2_55(G710,G4,G25);
  and AND2_56(G713,G4,G26);
  and AND2_57(G716,G4,G27);
  and AND2_58(G719,G4,G28);
  and AND2_59(G722,G4,G29);
  and AND2_60(G725,G4,G30);
  and AND2_61(G728,G4,G31);
  and AND2_62(G731,G4,G32);
  and AND2_63(G734,G5,G17);
  and AND2_64(G737,G5,G18);
  and AND2_65(G740,G5,G19);
  and AND2_66(G743,G5,G20);
  and AND2_67(G746,G5,G21);
  and AND2_68(G749,G5,G22);
  and AND2_69(G752,G5,G23);
  and AND2_70(G755,G5,G24);
  and AND2_71(G758,G5,G25);
  and AND2_72(G761,G5,G26);
  and AND2_73(G764,G5,G27);
  and AND2_74(G767,G5,G28);
  and AND2_75(G770,G5,G29);
  and AND2_76(G773,G5,G30);
  and AND2_77(G776,G5,G31);
  and AND2_78(G779,G5,G32);
  and AND2_79(G782,G6,G17);
  and AND2_80(G785,G6,G18);
  and AND2_81(G788,G6,G19);
  and AND2_82(G791,G6,G20);
  and AND2_83(G794,G6,G21);
  and AND2_84(G797,G6,G22);
  and AND2_85(G800,G6,G23);
  and AND2_86(G803,G6,G24);
  and AND2_87(G806,G6,G25);
  and AND2_88(G809,G6,G26);
  and AND2_89(G812,G6,G27);
  and AND2_90(G815,G6,G28);
  and AND2_91(G818,G6,G29);
  and AND2_92(G821,G6,G30);
  and AND2_93(G824,G6,G31);
  and AND2_94(G827,G6,G32);
  and AND2_95(G830,G7,G17);
  and AND2_96(G833,G7,G18);
  and AND2_97(G836,G7,G19);
  and AND2_98(G839,G7,G20);
  and AND2_99(G842,G7,G21);
  and AND2_100(G845,G7,G22);
  and AND2_101(G848,G7,G23);
  and AND2_102(G851,G7,G24);
  and AND2_103(G854,G7,G25);
  and AND2_104(G857,G7,G26);
  and AND2_105(G860,G7,G27);
  and AND2_106(G863,G7,G28);
  and AND2_107(G866,G7,G29);
  and AND2_108(G869,G7,G30);
  and AND2_109(G872,G7,G31);
  and AND2_110(G875,G7,G32);
  and AND2_111(G878,G8,G17);
  and AND2_112(G881,G8,G18);
  and AND2_113(G884,G8,G19);
  and AND2_114(G887,G8,G20);
  and AND2_115(G890,G8,G21);
  and AND2_116(G893,G8,G22);
  and AND2_117(G896,G8,G23);
  and AND2_118(G899,G8,G24);
  and AND2_119(G902,G8,G25);
  and AND2_120(G905,G8,G26);
  and AND2_121(G908,G8,G27);
  and AND2_122(G911,G8,G28);
  and AND2_123(G914,G8,G29);
  and AND2_124(G917,G8,G30);
  and AND2_125(G920,G8,G31);
  and AND2_126(G923,G8,G32);
  and AND2_127(G926,G9,G17);
  and AND2_128(G929,G9,G18);
  and AND2_129(G932,G9,G19);
  and AND2_130(G935,G9,G20);
  and AND2_131(G938,G9,G21);
  and AND2_132(G941,G9,G22);
  and AND2_133(G944,G9,G23);
  and AND2_134(G947,G9,G24);
  and AND2_135(G950,G9,G25);
  and AND2_136(G953,G9,G26);
  and AND2_137(G956,G9,G27);
  and AND2_138(G959,G9,G28);
  and AND2_139(G962,G9,G29);
  and AND2_140(G965,G9,G30);
  and AND2_141(G968,G9,G31);
  and AND2_142(G971,G9,G32);
  and AND2_143(G974,G10,G17);
  and AND2_144(G977,G10,G18);
  and AND2_145(G980,G10,G19);
  and AND2_146(G983,G10,G20);
  and AND2_147(G986,G10,G21);
  and AND2_148(G989,G10,G22);
  and AND2_149(G992,G10,G23);
  and AND2_150(G995,G10,G24);
  and AND2_151(G998,G10,G25);
  and AND2_152(G1001,G10,G26);
  and AND2_153(G1004,G10,G27);
  and AND2_154(G1007,G10,G28);
  and AND2_155(G1010,G10,G29);
  and AND2_156(G1013,G10,G30);
  and AND2_157(G1016,G10,G31);
  and AND2_158(G1019,G10,G32);
  and AND2_159(G1022,G11,G17);
  and AND2_160(G1025,G11,G18);
  and AND2_161(G1028,G11,G19);
  and AND2_162(G1031,G11,G20);
  and AND2_163(G1034,G11,G21);
  and AND2_164(G1037,G11,G22);
  and AND2_165(G1040,G11,G23);
  and AND2_166(G1043,G11,G24);
  and AND2_167(G1046,G11,G25);
  and AND2_168(G1049,G11,G26);
  and AND2_169(G1052,G11,G27);
  and AND2_170(G1055,G11,G28);
  and AND2_171(G1058,G11,G29);
  and AND2_172(G1061,G11,G30);
  and AND2_173(G1064,G11,G31);
  and AND2_174(G1067,G11,G32);
  and AND2_175(G1070,G12,G17);
  and AND2_176(G1073,G12,G18);
  and AND2_177(G1076,G12,G19);
  and AND2_178(G1079,G12,G20);
  and AND2_179(G1082,G12,G21);
  and AND2_180(G1085,G12,G22);
  and AND2_181(G1088,G12,G23);
  and AND2_182(G1091,G12,G24);
  and AND2_183(G1094,G12,G25);
  and AND2_184(G1097,G12,G26);
  and AND2_185(G1100,G12,G27);
  and AND2_186(G1103,G12,G28);
  and AND2_187(G1106,G12,G29);
  and AND2_188(G1109,G12,G30);
  and AND2_189(G1112,G12,G31);
  and AND2_190(G1115,G12,G32);
  and AND2_191(G1118,G13,G17);
  and AND2_192(G1121,G13,G18);
  and AND2_193(G1124,G13,G19);
  and AND2_194(G1127,G13,G20);
  and AND2_195(G1130,G13,G21);
  and AND2_196(G1133,G13,G22);
  and AND2_197(G1136,G13,G23);
  and AND2_198(G1139,G13,G24);
  and AND2_199(G1142,G13,G25);
  and AND2_200(G1145,G13,G26);
  and AND2_201(G1148,G13,G27);
  and AND2_202(G1151,G13,G28);
  and AND2_203(G1154,G13,G29);
  and AND2_204(G1157,G13,G30);
  and AND2_205(G1160,G13,G31);
  and AND2_206(G1163,G13,G32);
  and AND2_207(G1166,G14,G17);
  and AND2_208(G1169,G14,G18);
  and AND2_209(G1172,G14,G19);
  and AND2_210(G1175,G14,G20);
  and AND2_211(G1178,G14,G21);
  and AND2_212(G1181,G14,G22);
  and AND2_213(G1184,G14,G23);
  and AND2_214(G1187,G14,G24);
  and AND2_215(G1190,G14,G25);
  and AND2_216(G1193,G14,G26);
  and AND2_217(G1196,G14,G27);
  and AND2_218(G1199,G14,G28);
  and AND2_219(G1202,G14,G29);
  and AND2_220(G1205,G14,G30);
  and AND2_221(G1208,G14,G31);
  and AND2_222(G1211,G14,G32);
  and AND2_223(G1214,G15,G17);
  and AND2_224(G1217,G15,G18);
  and AND2_225(G1220,G15,G19);
  and AND2_226(G1223,G15,G20);
  and AND2_227(G1226,G15,G21);
  and AND2_228(G1229,G15,G22);
  and AND2_229(G1232,G15,G23);
  and AND2_230(G1235,G15,G24);
  and AND2_231(G1238,G15,G25);
  and AND2_232(G1241,G15,G26);
  and AND2_233(G1244,G15,G27);
  and AND2_234(G1247,G15,G28);
  and AND2_235(G1250,G15,G29);
  and AND2_236(G1253,G15,G30);
  and AND2_237(G1256,G15,G31);
  and AND2_238(G1259,G15,G32);
  and AND2_239(G1262,G16,G17);
  and AND2_240(G1265,G16,G18);
  and AND2_241(G1268,G16,G19);
  and AND2_242(G1271,G16,G20);
  and AND2_243(G1274,G16,G21);
  and AND2_244(G1277,G16,G22);
  and AND2_245(G1280,G16,G23);
  and AND2_246(G1283,G16,G24);
  and AND2_247(G1286,G16,G25);
  and AND2_248(G1289,G16,G26);
  and AND2_249(G1292,G16,G27);
  and AND2_250(G1295,G16,G28);
  and AND2_251(G1298,G16,G29);
  and AND2_252(G1301,G16,G30);
  and AND2_253(G1304,G16,G31);
  and AND2_254(G1307,G16,G32);
  not NOT_0(G1310,G590);
  not NOT_1(G1314,G638);
  not NOT_2(G1318,G686);
  not NOT_3(G1322,G734);
  not NOT_4(G1326,G782);
  not NOT_5(G1330,G830);
  not NOT_6(G1334,G878);
  not NOT_7(G1338,G926);
  not NOT_8(G1342,G974);
  not NOT_9(G1346,G1022);
  not NOT_10(G1350,G1070);
  not NOT_11(G1354,G1118);
  not NOT_12(G1358,G1166);
  not NOT_13(G1362,G1214);
  not NOT_14(G1366,G1262);
  nor NOR2_0(G1370,G590,G1310);
  not NOT_15(G1371,G1310);
  nor NOR2_1(G1372,G638,G1314);
  not NOT_16(G1373,G1314);
  nor NOR2_2(G1374,G686,G1318);
  not NOT_17(G1375,G1318);
  nor NOR2_3(G1376,G734,G1322);
  not NOT_18(G1377,G1322);
  nor NOR2_4(G1378,G782,G1326);
  not NOT_19(G1379,G1326);
  nor NOR2_5(G1380,G830,G1330);
  not NOT_20(G1381,G1330);
  nor NOR2_6(G1382,G878,G1334);
  not NOT_21(G1383,G1334);
  nor NOR2_7(G1384,G926,G1338);
  not NOT_22(G1385,G1338);
  nor NOR2_8(G1386,G974,G1342);
  not NOT_23(G1387,G1342);
  nor NOR2_9(G1388,G1022,G1346);
  not NOT_24(G1389,G1346);
  nor NOR2_10(G1390,G1070,G1350);
  not NOT_25(G1391,G1350);
  nor NOR2_11(G1392,G1118,G1354);
  not NOT_26(G1393,G1354);
  nor NOR2_12(G1394,G1166,G1358);
  not NOT_27(G1395,G1358);
  nor NOR2_13(G1396,G1214,G1362);
  not NOT_28(G1397,G1362);
  nor NOR2_14(G1398,G1262,G1366);
  not NOT_29(G1399,G1366);
  nor NOR2_15(G1400,G1370,G1371);
  nor NOR2_16(G1403,G1372,G1373);
  nor NOR2_17(G1406,G1374,G1375);
  nor NOR2_18(G1409,G1376,G1377);
  nor NOR2_19(G1412,G1378,G1379);
  nor NOR2_20(G1415,G1380,G1381);
  nor NOR2_21(G1418,G1382,G1383);
  nor NOR2_22(G1421,G1384,G1385);
  nor NOR2_23(G1424,G1386,G1387);
  nor NOR2_24(G1427,G1388,G1389);
  nor NOR2_25(G1430,G1390,G1391);
  nor NOR2_26(G1433,G1392,G1393);
  nor NOR2_27(G1436,G1394,G1395);
  nor NOR2_28(G1439,G1396,G1397);
  nor NOR2_29(G1442,G1398,G1399);
  nor NOR2_30(G1445,G1400,G545);
  nor NOR2_31(G1449,G1403,G593);
  nor NOR2_32(G1453,G1406,G641);
  nor NOR2_33(G1457,G1409,G689);
  nor NOR2_34(G1461,G1412,G737);
  nor NOR2_35(G1465,G1415,G785);
  nor NOR2_36(G1469,G1418,G833);
  nor NOR2_37(G1473,G1421,G881);
  nor NOR2_38(G1477,G1424,G929);
  nor NOR2_39(G1481,G1427,G977);
  nor NOR2_40(G1485,G1430,G1025);
  nor NOR2_41(G1489,G1433,G1073);
  nor NOR2_42(G1493,G1436,G1121);
  nor NOR2_43(G1497,G1439,G1169);
  nor NOR2_44(G1501,G1442,G1217);
  nor NOR2_45(G1505,G1400,G1445);
  nor NOR2_46(G1506,G1445,G545);
  nor NOR2_47(G1507,G1310,G1445);
  nor NOR2_48(G1510,G1403,G1449);
  nor NOR2_49(G1511,G1449,G593);
  nor NOR2_50(G1512,G1314,G1449);
  nor NOR2_51(G1515,G1406,G1453);
  nor NOR2_52(G1516,G1453,G641);
  nor NOR2_53(G1517,G1318,G1453);
  nor NOR2_54(G1520,G1409,G1457);
  nor NOR2_55(G1521,G1457,G689);
  nor NOR2_56(G1522,G1322,G1457);
  nor NOR2_57(G1525,G1412,G1461);
  nor NOR2_58(G1526,G1461,G737);
  nor NOR2_59(G1527,G1326,G1461);
  nor NOR2_60(G1530,G1415,G1465);
  nor NOR2_61(G1531,G1465,G785);
  nor NOR2_62(G1532,G1330,G1465);
  nor NOR2_63(G1535,G1418,G1469);
  nor NOR2_64(G1536,G1469,G833);
  nor NOR2_65(G1537,G1334,G1469);
  nor NOR2_66(G1540,G1421,G1473);
  nor NOR2_67(G1541,G1473,G881);
  nor NOR2_68(G1542,G1338,G1473);
  nor NOR2_69(G1545,G1424,G1477);
  nor NOR2_70(G1546,G1477,G929);
  nor NOR2_71(G1547,G1342,G1477);
  nor NOR2_72(G1550,G1427,G1481);
  nor NOR2_73(G1551,G1481,G977);
  nor NOR2_74(G1552,G1346,G1481);
  nor NOR2_75(G1555,G1430,G1485);
  nor NOR2_76(G1556,G1485,G1025);
  nor NOR2_77(G1557,G1350,G1485);
  nor NOR2_78(G1560,G1433,G1489);
  nor NOR2_79(G1561,G1489,G1073);
  nor NOR2_80(G1562,G1354,G1489);
  nor NOR2_81(G1565,G1436,G1493);
  nor NOR2_82(G1566,G1493,G1121);
  nor NOR2_83(G1567,G1358,G1493);
  nor NOR2_84(G1570,G1439,G1497);
  nor NOR2_85(G1571,G1497,G1169);
  nor NOR2_86(G1572,G1362,G1497);
  nor NOR2_87(G1575,G1442,G1501);
  nor NOR2_88(G1576,G1501,G1217);
  nor NOR2_89(G1577,G1366,G1501);
  nor NOR2_90(G1580,G1510,G1511);
  nor NOR2_91(G1583,G1515,G1516);
  nor NOR2_92(G1586,G1520,G1521);
  nor NOR2_93(G1589,G1525,G1526);
  nor NOR2_94(G1592,G1530,G1531);
  nor NOR2_95(G1595,G1535,G1536);
  nor NOR2_96(G1598,G1540,G1541);
  nor NOR2_97(G1601,G1545,G1546);
  nor NOR2_98(G1604,G1550,G1551);
  nor NOR2_99(G1607,G1555,G1556);
  nor NOR2_100(G1610,G1560,G1561);
  nor NOR2_101(G1613,G1565,G1566);
  nor NOR2_102(G1616,G1570,G1571);
  nor NOR2_103(G1619,G1575,G1576);
  nor NOR2_104(G1622,G1265,G1577);
  nor NOR2_105(G1626,G1580,G1507);
  nor NOR2_106(G1630,G1583,G1512);
  nor NOR2_107(G1634,G1586,G1517);
  nor NOR2_108(G1638,G1589,G1522);
  nor NOR2_109(G1642,G1592,G1527);
  nor NOR2_110(G1646,G1595,G1532);
  nor NOR2_111(G1650,G1598,G1537);
  nor NOR2_112(G1654,G1601,G1542);
  nor NOR2_113(G1658,G1604,G1547);
  nor NOR2_114(G1662,G1607,G1552);
  nor NOR2_115(G1666,G1610,G1557);
  nor NOR2_116(G1670,G1613,G1562);
  nor NOR2_117(G1674,G1616,G1567);
  nor NOR2_118(G1678,G1619,G1572);
  nor NOR2_119(G1682,G1265,G1622);
  nor NOR2_120(G1683,G1622,G1577);
  nor NOR2_121(G1684,G1580,G1626);
  nor NOR2_122(G1685,G1626,G1507);
  nor NOR2_123(G1686,G1583,G1630);
  nor NOR2_124(G1687,G1630,G1512);
  nor NOR2_125(G1688,G1586,G1634);
  nor NOR2_126(G1689,G1634,G1517);
  nor NOR2_127(G1690,G1589,G1638);
  nor NOR2_128(G1691,G1638,G1522);
  nor NOR2_129(G1692,G1592,G1642);
  nor NOR2_130(G1693,G1642,G1527);
  nor NOR2_131(G1694,G1595,G1646);
  nor NOR2_132(G1695,G1646,G1532);
  nor NOR2_133(G1696,G1598,G1650);
  nor NOR2_134(G1697,G1650,G1537);
  nor NOR2_135(G1698,G1601,G1654);
  nor NOR2_136(G1699,G1654,G1542);
  nor NOR2_137(G1700,G1604,G1658);
  nor NOR2_138(G1701,G1658,G1547);
  nor NOR2_139(G1702,G1607,G1662);
  nor NOR2_140(G1703,G1662,G1552);
  nor NOR2_141(G1704,G1610,G1666);
  nor NOR2_142(G1705,G1666,G1557);
  nor NOR2_143(G1706,G1613,G1670);
  nor NOR2_144(G1707,G1670,G1562);
  nor NOR2_145(G1708,G1616,G1674);
  nor NOR2_146(G1709,G1674,G1567);
  nor NOR2_147(G1710,G1619,G1678);
  nor NOR2_148(G1711,G1678,G1572);
  nor NOR2_149(G1712,G1682,G1683);
  nor NOR2_150(G1715,G1684,G1685);
  nor NOR2_151(G1718,G1686,G1687);
  nor NOR2_152(G1721,G1688,G1689);
  nor NOR2_153(G1724,G1690,G1691);
  nor NOR2_154(G1727,G1692,G1693);
  nor NOR2_155(G1730,G1694,G1695);
  nor NOR2_156(G1733,G1696,G1697);
  nor NOR2_157(G1736,G1698,G1699);
  nor NOR2_158(G1739,G1700,G1701);
  nor NOR2_159(G1742,G1702,G1703);
  nor NOR2_160(G1745,G1704,G1705);
  nor NOR2_161(G1748,G1706,G1707);
  nor NOR2_162(G1751,G1708,G1709);
  nor NOR2_163(G1754,G1710,G1711);
  nor NOR2_164(G1757,G1712,G1220);
  nor NOR2_165(G1761,G1715,G548);
  nor NOR2_166(G1765,G1718,G596);
  nor NOR2_167(G1769,G1721,G644);
  nor NOR2_168(G1773,G1724,G692);
  nor NOR2_169(G1777,G1727,G740);
  nor NOR2_170(G1781,G1730,G788);
  nor NOR2_171(G1785,G1733,G836);
  nor NOR2_172(G1789,G1736,G884);
  nor NOR2_173(G1793,G1739,G932);
  nor NOR2_174(G1797,G1742,G980);
  nor NOR2_175(G1801,G1745,G1028);
  nor NOR2_176(G1805,G1748,G1076);
  nor NOR2_177(G1809,G1751,G1124);
  nor NOR2_178(G1813,G1754,G1172);
  nor NOR2_179(G1817,G1712,G1757);
  nor NOR2_180(G1818,G1757,G1220);
  nor NOR2_181(G1819,G1622,G1757);
  nor NOR2_182(G1822,G1715,G1761);
  nor NOR2_183(G1823,G1761,G548);
  nor NOR2_184(G1824,G1626,G1761);
  nor NOR2_185(G1827,G1718,G1765);
  nor NOR2_186(G1828,G1765,G596);
  nor NOR2_187(G1829,G1630,G1765);
  nor NOR2_188(G1832,G1721,G1769);
  nor NOR2_189(G1833,G1769,G644);
  nor NOR2_190(G1834,G1634,G1769);
  nor NOR2_191(G1837,G1724,G1773);
  nor NOR2_192(G1838,G1773,G692);
  nor NOR2_193(G1839,G1638,G1773);
  nor NOR2_194(G1842,G1727,G1777);
  nor NOR2_195(G1843,G1777,G740);
  nor NOR2_196(G1844,G1642,G1777);
  nor NOR2_197(G1847,G1730,G1781);
  nor NOR2_198(G1848,G1781,G788);
  nor NOR2_199(G1849,G1646,G1781);
  nor NOR2_200(G1852,G1733,G1785);
  nor NOR2_201(G1853,G1785,G836);
  nor NOR2_202(G1854,G1650,G1785);
  nor NOR2_203(G1857,G1736,G1789);
  nor NOR2_204(G1858,G1789,G884);
  nor NOR2_205(G1859,G1654,G1789);
  nor NOR2_206(G1862,G1739,G1793);
  nor NOR2_207(G1863,G1793,G932);
  nor NOR2_208(G1864,G1658,G1793);
  nor NOR2_209(G1867,G1742,G1797);
  nor NOR2_210(G1868,G1797,G980);
  nor NOR2_211(G1869,G1662,G1797);
  nor NOR2_212(G1872,G1745,G1801);
  nor NOR2_213(G1873,G1801,G1028);
  nor NOR2_214(G1874,G1666,G1801);
  nor NOR2_215(G1877,G1748,G1805);
  nor NOR2_216(G1878,G1805,G1076);
  nor NOR2_217(G1879,G1670,G1805);
  nor NOR2_218(G1882,G1751,G1809);
  nor NOR2_219(G1883,G1809,G1124);
  nor NOR2_220(G1884,G1674,G1809);
  nor NOR2_221(G1887,G1754,G1813);
  nor NOR2_222(G1888,G1813,G1172);
  nor NOR2_223(G1889,G1678,G1813);
  nor NOR2_224(G1892,G1817,G1818);
  nor NOR2_225(G1895,G1268,G1819);
  nor NOR2_226(G1899,G1827,G1828);
  nor NOR2_227(G1902,G1832,G1833);
  nor NOR2_228(G1905,G1837,G1838);
  nor NOR2_229(G1908,G1842,G1843);
  nor NOR2_230(G1911,G1847,G1848);
  nor NOR2_231(G1914,G1852,G1853);
  nor NOR2_232(G1917,G1857,G1858);
  nor NOR2_233(G1920,G1862,G1863);
  nor NOR2_234(G1923,G1867,G1868);
  nor NOR2_235(G1926,G1872,G1873);
  nor NOR2_236(G1929,G1877,G1878);
  nor NOR2_237(G1932,G1882,G1883);
  nor NOR2_238(G1935,G1887,G1888);
  nor NOR2_239(G1938,G1892,G1889);
  nor NOR2_240(G1942,G1268,G1895);
  nor NOR2_241(G1943,G1895,G1819);
  nor NOR2_242(G1944,G1899,G1824);
  nor NOR2_243(G1948,G1902,G1829);
  nor NOR2_244(G1952,G1905,G1834);
  nor NOR2_245(G1956,G1908,G1839);
  nor NOR2_246(G1960,G1911,G1844);
  nor NOR2_247(G1964,G1914,G1849);
  nor NOR2_248(G1968,G1917,G1854);
  nor NOR2_249(G1972,G1920,G1859);
  nor NOR2_250(G1976,G1923,G1864);
  nor NOR2_251(G1980,G1926,G1869);
  nor NOR2_252(G1984,G1929,G1874);
  nor NOR2_253(G1988,G1932,G1879);
  nor NOR2_254(G1992,G1935,G1884);
  nor NOR2_255(G1996,G1892,G1938);
  nor NOR2_256(G1997,G1938,G1889);
  nor NOR2_257(G1998,G1942,G1943);
  nor NOR2_258(G2001,G1899,G1944);
  nor NOR2_259(G2002,G1944,G1824);
  nor NOR2_260(G2003,G1902,G1948);
  nor NOR2_261(G2004,G1948,G1829);
  nor NOR2_262(G2005,G1905,G1952);
  nor NOR2_263(G2006,G1952,G1834);
  nor NOR2_264(G2007,G1908,G1956);
  nor NOR2_265(G2008,G1956,G1839);
  nor NOR2_266(G2009,G1911,G1960);
  nor NOR2_267(G2010,G1960,G1844);
  nor NOR2_268(G2011,G1914,G1964);
  nor NOR2_269(G2012,G1964,G1849);
  nor NOR2_270(G2013,G1917,G1968);
  nor NOR2_271(G2014,G1968,G1854);
  nor NOR2_272(G2015,G1920,G1972);
  nor NOR2_273(G2016,G1972,G1859);
  nor NOR2_274(G2017,G1923,G1976);
  nor NOR2_275(G2018,G1976,G1864);
  nor NOR2_276(G2019,G1926,G1980);
  nor NOR2_277(G2020,G1980,G1869);
  nor NOR2_278(G2021,G1929,G1984);
  nor NOR2_279(G2022,G1984,G1874);
  nor NOR2_280(G2023,G1932,G1988);
  nor NOR2_281(G2024,G1988,G1879);
  nor NOR2_282(G2025,G1935,G1992);
  nor NOR2_283(G2026,G1992,G1884);
  nor NOR2_284(G2027,G1996,G1997);
  nor NOR2_285(G2030,G1998,G1223);
  nor NOR2_286(G2034,G2001,G2002);
  nor NOR2_287(G2037,G2003,G2004);
  nor NOR2_288(G2040,G2005,G2006);
  nor NOR2_289(G2043,G2007,G2008);
  nor NOR2_290(G2046,G2009,G2010);
  nor NOR2_291(G2049,G2011,G2012);
  nor NOR2_292(G2052,G2013,G2014);
  nor NOR2_293(G2055,G2015,G2016);
  nor NOR2_294(G2058,G2017,G2018);
  nor NOR2_295(G2061,G2019,G2020);
  nor NOR2_296(G2064,G2021,G2022);
  nor NOR2_297(G2067,G2023,G2024);
  nor NOR2_298(G2070,G2025,G2026);
  nor NOR2_299(G2073,G2027,G1175);
  nor NOR2_300(G2077,G1998,G2030);
  nor NOR2_301(G2078,G2030,G1223);
  nor NOR2_302(G2079,G1895,G2030);
  nor NOR2_303(G2082,G2034,G551);
  nor NOR2_304(G2086,G2037,G599);
  nor NOR2_305(G2090,G2040,G647);
  nor NOR2_306(G2094,G2043,G695);
  nor NOR2_307(G2098,G2046,G743);
  nor NOR2_308(G2102,G2049,G791);
  nor NOR2_309(G2106,G2052,G839);
  nor NOR2_310(G2110,G2055,G887);
  nor NOR2_311(G2114,G2058,G935);
  nor NOR2_312(G2118,G2061,G983);
  nor NOR2_313(G2122,G2064,G1031);
  nor NOR2_314(G2126,G2067,G1079);
  nor NOR2_315(G2130,G2070,G1127);
  nor NOR2_316(G2134,G2027,G2073);
  nor NOR2_317(G2135,G2073,G1175);
  nor NOR2_318(G2136,G1938,G2073);
  nor NOR2_319(G2139,G2077,G2078);
  nor NOR2_320(G2142,G1271,G2079);
  nor NOR2_321(G2146,G2034,G2082);
  nor NOR2_322(G2147,G2082,G551);
  nor NOR2_323(G2148,G1944,G2082);
  nor NOR2_324(G2151,G2037,G2086);
  nor NOR2_325(G2152,G2086,G599);
  nor NOR2_326(G2153,G1948,G2086);
  nor NOR2_327(G2156,G2040,G2090);
  nor NOR2_328(G2157,G2090,G647);
  nor NOR2_329(G2158,G1952,G2090);
  nor NOR2_330(G2161,G2043,G2094);
  nor NOR2_331(G2162,G2094,G695);
  nor NOR2_332(G2163,G1956,G2094);
  nor NOR2_333(G2166,G2046,G2098);
  nor NOR2_334(G2167,G2098,G743);
  nor NOR2_335(G2168,G1960,G2098);
  nor NOR2_336(G2171,G2049,G2102);
  nor NOR2_337(G2172,G2102,G791);
  nor NOR2_338(G2173,G1964,G2102);
  nor NOR2_339(G2176,G2052,G2106);
  nor NOR2_340(G2177,G2106,G839);
  nor NOR2_341(G2178,G1968,G2106);
  nor NOR2_342(G2181,G2055,G2110);
  nor NOR2_343(G2182,G2110,G887);
  nor NOR2_344(G2183,G1972,G2110);
  nor NOR2_345(G2186,G2058,G2114);
  nor NOR2_346(G2187,G2114,G935);
  nor NOR2_347(G2188,G1976,G2114);
  nor NOR2_348(G2191,G2061,G2118);
  nor NOR2_349(G2192,G2118,G983);
  nor NOR2_350(G2193,G1980,G2118);
  nor NOR2_351(G2196,G2064,G2122);
  nor NOR2_352(G2197,G2122,G1031);
  nor NOR2_353(G2198,G1984,G2122);
  nor NOR2_354(G2201,G2067,G2126);
  nor NOR2_355(G2202,G2126,G1079);
  nor NOR2_356(G2203,G1988,G2126);
  nor NOR2_357(G2206,G2070,G2130);
  nor NOR2_358(G2207,G2130,G1127);
  nor NOR2_359(G2208,G1992,G2130);
  nor NOR2_360(G2211,G2134,G2135);
  nor NOR2_361(G2214,G2139,G2136);
  nor NOR2_362(G2218,G1271,G2142);
  nor NOR2_363(G2219,G2142,G2079);
  nor NOR2_364(G2220,G2151,G2152);
  nor NOR2_365(G2223,G2156,G2157);
  nor NOR2_366(G2226,G2161,G2162);
  nor NOR2_367(G2229,G2166,G2167);
  nor NOR2_368(G2232,G2171,G2172);
  nor NOR2_369(G2235,G2176,G2177);
  nor NOR2_370(G2238,G2181,G2182);
  nor NOR2_371(G2241,G2186,G2187);
  nor NOR2_372(G2244,G2191,G2192);
  nor NOR2_373(G2247,G2196,G2197);
  nor NOR2_374(G2250,G2201,G2202);
  nor NOR2_375(G2253,G2206,G2207);
  nor NOR2_376(G2256,G2211,G2208);
  nor NOR2_377(G2260,G2139,G2214);
  nor NOR2_378(G2261,G2214,G2136);
  nor NOR2_379(G2262,G2218,G2219);
  nor NOR2_380(G2265,G2220,G2148);
  nor NOR2_381(G2269,G2223,G2153);
  nor NOR2_382(G2273,G2226,G2158);
  nor NOR2_383(G2277,G2229,G2163);
  nor NOR2_384(G2281,G2232,G2168);
  nor NOR2_385(G2285,G2235,G2173);
  nor NOR2_386(G2289,G2238,G2178);
  nor NOR2_387(G2293,G2241,G2183);
  nor NOR2_388(G2297,G2244,G2188);
  nor NOR2_389(G2301,G2247,G2193);
  nor NOR2_390(G2305,G2250,G2198);
  nor NOR2_391(G2309,G2253,G2203);
  nor NOR2_392(G2313,G2211,G2256);
  nor NOR2_393(G2314,G2256,G2208);
  nor NOR2_394(G2315,G2260,G2261);
  nor NOR2_395(G2318,G2262,G1226);
  nor NOR2_396(G2322,G2220,G2265);
  nor NOR2_397(G2323,G2265,G2148);
  nor NOR2_398(G2324,G2223,G2269);
  nor NOR2_399(G2325,G2269,G2153);
  nor NOR2_400(G2326,G2226,G2273);
  nor NOR2_401(G2327,G2273,G2158);
  nor NOR2_402(G2328,G2229,G2277);
  nor NOR2_403(G2329,G2277,G2163);
  nor NOR2_404(G2330,G2232,G2281);
  nor NOR2_405(G2331,G2281,G2168);
  nor NOR2_406(G2332,G2235,G2285);
  nor NOR2_407(G2333,G2285,G2173);
  nor NOR2_408(G2334,G2238,G2289);
  nor NOR2_409(G2335,G2289,G2178);
  nor NOR2_410(G2336,G2241,G2293);
  nor NOR2_411(G2337,G2293,G2183);
  nor NOR2_412(G2338,G2244,G2297);
  nor NOR2_413(G2339,G2297,G2188);
  nor NOR2_414(G2340,G2247,G2301);
  nor NOR2_415(G2341,G2301,G2193);
  nor NOR2_416(G2342,G2250,G2305);
  nor NOR2_417(G2343,G2305,G2198);
  nor NOR2_418(G2344,G2253,G2309);
  nor NOR2_419(G2345,G2309,G2203);
  nor NOR2_420(G2346,G2313,G2314);
  nor NOR2_421(G2349,G2315,G1178);
  nor NOR2_422(G2353,G2262,G2318);
  nor NOR2_423(G2354,G2318,G1226);
  nor NOR2_424(G2355,G2142,G2318);
  nor NOR2_425(G2358,G2322,G2323);
  nor NOR2_426(G2361,G2324,G2325);
  nor NOR2_427(G2364,G2326,G2327);
  nor NOR2_428(G2367,G2328,G2329);
  nor NOR2_429(G2370,G2330,G2331);
  nor NOR2_430(G2373,G2332,G2333);
  nor NOR2_431(G2376,G2334,G2335);
  nor NOR2_432(G2379,G2336,G2337);
  nor NOR2_433(G2382,G2338,G2339);
  nor NOR2_434(G2385,G2340,G2341);
  nor NOR2_435(G2388,G2342,G2343);
  nor NOR2_436(G2391,G2344,G2345);
  nor NOR2_437(G2394,G2346,G1130);
  nor NOR2_438(G2398,G2315,G2349);
  nor NOR2_439(G2399,G2349,G1178);
  nor NOR2_440(G2400,G2214,G2349);
  nor NOR2_441(G2403,G2353,G2354);
  nor NOR2_442(G2406,G1274,G2355);
  nor NOR2_443(G2410,G2358,G554);
  nor NOR2_444(G2414,G2361,G602);
  nor NOR2_445(G2418,G2364,G650);
  nor NOR2_446(G2422,G2367,G698);
  nor NOR2_447(G2426,G2370,G746);
  nor NOR2_448(G2430,G2373,G794);
  nor NOR2_449(G2434,G2376,G842);
  nor NOR2_450(G2438,G2379,G890);
  nor NOR2_451(G2442,G2382,G938);
  nor NOR2_452(G2446,G2385,G986);
  nor NOR2_453(G2450,G2388,G1034);
  nor NOR2_454(G2454,G2391,G1082);
  nor NOR2_455(G2458,G2346,G2394);
  nor NOR2_456(G2459,G2394,G1130);
  nor NOR2_457(G2460,G2256,G2394);
  nor NOR2_458(G2463,G2398,G2399);
  nor NOR2_459(G2466,G2403,G2400);
  nor NOR2_460(G2470,G1274,G2406);
  nor NOR2_461(G2471,G2406,G2355);
  nor NOR2_462(G2472,G2358,G2410);
  nor NOR2_463(G2473,G2410,G554);
  nor NOR2_464(G2474,G2265,G2410);
  nor NOR2_465(G2477,G2361,G2414);
  nor NOR2_466(G2478,G2414,G602);
  nor NOR2_467(G2479,G2269,G2414);
  nor NOR2_468(G2482,G2364,G2418);
  nor NOR2_469(G2483,G2418,G650);
  nor NOR2_470(G2484,G2273,G2418);
  nor NOR2_471(G2487,G2367,G2422);
  nor NOR2_472(G2488,G2422,G698);
  nor NOR2_473(G2489,G2277,G2422);
  nor NOR2_474(G2492,G2370,G2426);
  nor NOR2_475(G2493,G2426,G746);
  nor NOR2_476(G2494,G2281,G2426);
  nor NOR2_477(G2497,G2373,G2430);
  nor NOR2_478(G2498,G2430,G794);
  nor NOR2_479(G2499,G2285,G2430);
  nor NOR2_480(G2502,G2376,G2434);
  nor NOR2_481(G2503,G2434,G842);
  nor NOR2_482(G2504,G2289,G2434);
  nor NOR2_483(G2507,G2379,G2438);
  nor NOR2_484(G2508,G2438,G890);
  nor NOR2_485(G2509,G2293,G2438);
  nor NOR2_486(G2512,G2382,G2442);
  nor NOR2_487(G2513,G2442,G938);
  nor NOR2_488(G2514,G2297,G2442);
  nor NOR2_489(G2517,G2385,G2446);
  nor NOR2_490(G2518,G2446,G986);
  nor NOR2_491(G2519,G2301,G2446);
  nor NOR2_492(G2522,G2388,G2450);
  nor NOR2_493(G2523,G2450,G1034);
  nor NOR2_494(G2524,G2305,G2450);
  nor NOR2_495(G2527,G2391,G2454);
  nor NOR2_496(G2528,G2454,G1082);
  nor NOR2_497(G2529,G2309,G2454);
  nor NOR2_498(G2532,G2458,G2459);
  nor NOR2_499(G2535,G2463,G2460);
  nor NOR2_500(G2539,G2403,G2466);
  nor NOR2_501(G2540,G2466,G2400);
  nor NOR2_502(G2541,G2470,G2471);
  nor NOR2_503(G2544,G2477,G2478);
  nor NOR2_504(G2547,G2482,G2483);
  nor NOR2_505(G2550,G2487,G2488);
  nor NOR2_506(G2553,G2492,G2493);
  nor NOR2_507(G2556,G2497,G2498);
  nor NOR2_508(G2559,G2502,G2503);
  nor NOR2_509(G2562,G2507,G2508);
  nor NOR2_510(G2565,G2512,G2513);
  nor NOR2_511(G2568,G2517,G2518);
  nor NOR2_512(G2571,G2522,G2523);
  nor NOR2_513(G2574,G2527,G2528);
  nor NOR2_514(G2577,G2532,G2529);
  nor NOR2_515(G2581,G2463,G2535);
  nor NOR2_516(G2582,G2535,G2460);
  nor NOR2_517(G2583,G2539,G2540);
  nor NOR2_518(G2586,G2541,G1229);
  nor NOR2_519(G2590,G2544,G2474);
  nor NOR2_520(G2594,G2547,G2479);
  nor NOR2_521(G2598,G2550,G2484);
  nor NOR2_522(G2602,G2553,G2489);
  nor NOR2_523(G2606,G2556,G2494);
  nor NOR2_524(G2610,G2559,G2499);
  nor NOR2_525(G2614,G2562,G2504);
  nor NOR2_526(G2618,G2565,G2509);
  nor NOR2_527(G2622,G2568,G2514);
  nor NOR2_528(G2626,G2571,G2519);
  nor NOR2_529(G2630,G2574,G2524);
  nor NOR2_530(G2634,G2532,G2577);
  nor NOR2_531(G2635,G2577,G2529);
  nor NOR2_532(G2636,G2581,G2582);
  nor NOR2_533(G2639,G2583,G1181);
  nor NOR2_534(G2643,G2541,G2586);
  nor NOR2_535(G2644,G2586,G1229);
  nor NOR2_536(G2645,G2406,G2586);
  nor NOR2_537(G2648,G2544,G2590);
  nor NOR2_538(G2649,G2590,G2474);
  nor NOR2_539(G2650,G2547,G2594);
  nor NOR2_540(G2651,G2594,G2479);
  nor NOR2_541(G2652,G2550,G2598);
  nor NOR2_542(G2653,G2598,G2484);
  nor NOR2_543(G2654,G2553,G2602);
  nor NOR2_544(G2655,G2602,G2489);
  nor NOR2_545(G2656,G2556,G2606);
  nor NOR2_546(G2657,G2606,G2494);
  nor NOR2_547(G2658,G2559,G2610);
  nor NOR2_548(G2659,G2610,G2499);
  nor NOR2_549(G2660,G2562,G2614);
  nor NOR2_550(G2661,G2614,G2504);
  nor NOR2_551(G2662,G2565,G2618);
  nor NOR2_552(G2663,G2618,G2509);
  nor NOR2_553(G2664,G2568,G2622);
  nor NOR2_554(G2665,G2622,G2514);
  nor NOR2_555(G2666,G2571,G2626);
  nor NOR2_556(G2667,G2626,G2519);
  nor NOR2_557(G2668,G2574,G2630);
  nor NOR2_558(G2669,G2630,G2524);
  nor NOR2_559(G2670,G2634,G2635);
  nor NOR2_560(G2673,G2636,G1133);
  nor NOR2_561(G2677,G2583,G2639);
  nor NOR2_562(G2678,G2639,G1181);
  nor NOR2_563(G2679,G2466,G2639);
  nor NOR2_564(G2682,G2643,G2644);
  nor NOR2_565(G2685,G1277,G2645);
  nor NOR2_566(G2689,G2648,G2649);
  nor NOR2_567(G2692,G2650,G2651);
  nor NOR2_568(G2695,G2652,G2653);
  nor NOR2_569(G2698,G2654,G2655);
  nor NOR2_570(G2701,G2656,G2657);
  nor NOR2_571(G2704,G2658,G2659);
  nor NOR2_572(G2707,G2660,G2661);
  nor NOR2_573(G2710,G2662,G2663);
  nor NOR2_574(G2713,G2664,G2665);
  nor NOR2_575(G2716,G2666,G2667);
  nor NOR2_576(G2719,G2668,G2669);
  nor NOR2_577(G2722,G2670,G1085);
  nor NOR2_578(G2726,G2636,G2673);
  nor NOR2_579(G2727,G2673,G1133);
  nor NOR2_580(G2728,G2535,G2673);
  nor NOR2_581(G2731,G2677,G2678);
  nor NOR2_582(G2734,G2682,G2679);
  nor NOR2_583(G2738,G1277,G2685);
  nor NOR2_584(G2739,G2685,G2645);
  nor NOR2_585(G2740,G2689,G557);
  nor NOR2_586(G2744,G2692,G605);
  nor NOR2_587(G2748,G2695,G653);
  nor NOR2_588(G2752,G2698,G701);
  nor NOR2_589(G2756,G2701,G749);
  nor NOR2_590(G2760,G2704,G797);
  nor NOR2_591(G2764,G2707,G845);
  nor NOR2_592(G2768,G2710,G893);
  nor NOR2_593(G2772,G2713,G941);
  nor NOR2_594(G2776,G2716,G989);
  nor NOR2_595(G2780,G2719,G1037);
  nor NOR2_596(G2784,G2670,G2722);
  nor NOR2_597(G2785,G2722,G1085);
  nor NOR2_598(G2786,G2577,G2722);
  nor NOR2_599(G2789,G2726,G2727);
  nor NOR2_600(G2792,G2731,G2728);
  nor NOR2_601(G2796,G2682,G2734);
  nor NOR2_602(G2797,G2734,G2679);
  nor NOR2_603(G2798,G2738,G2739);
  nor NOR2_604(G2801,G2689,G2740);
  nor NOR2_605(G2802,G2740,G557);
  nor NOR2_606(G2803,G2590,G2740);
  nor NOR2_607(G2806,G2692,G2744);
  nor NOR2_608(G2807,G2744,G605);
  nor NOR2_609(G2808,G2594,G2744);
  nor NOR2_610(G2811,G2695,G2748);
  nor NOR2_611(G2812,G2748,G653);
  nor NOR2_612(G2813,G2598,G2748);
  nor NOR2_613(G2816,G2698,G2752);
  nor NOR2_614(G2817,G2752,G701);
  nor NOR2_615(G2818,G2602,G2752);
  nor NOR2_616(G2821,G2701,G2756);
  nor NOR2_617(G2822,G2756,G749);
  nor NOR2_618(G2823,G2606,G2756);
  nor NOR2_619(G2826,G2704,G2760);
  nor NOR2_620(G2827,G2760,G797);
  nor NOR2_621(G2828,G2610,G2760);
  nor NOR2_622(G2831,G2707,G2764);
  nor NOR2_623(G2832,G2764,G845);
  nor NOR2_624(G2833,G2614,G2764);
  nor NOR2_625(G2836,G2710,G2768);
  nor NOR2_626(G2837,G2768,G893);
  nor NOR2_627(G2838,G2618,G2768);
  nor NOR2_628(G2841,G2713,G2772);
  nor NOR2_629(G2842,G2772,G941);
  nor NOR2_630(G2843,G2622,G2772);
  nor NOR2_631(G2846,G2716,G2776);
  nor NOR2_632(G2847,G2776,G989);
  nor NOR2_633(G2848,G2626,G2776);
  nor NOR2_634(G2851,G2719,G2780);
  nor NOR2_635(G2852,G2780,G1037);
  nor NOR2_636(G2853,G2630,G2780);
  nor NOR2_637(G2856,G2784,G2785);
  nor NOR2_638(G2859,G2789,G2786);
  nor NOR2_639(G2863,G2731,G2792);
  nor NOR2_640(G2864,G2792,G2728);
  nor NOR2_641(G2865,G2796,G2797);
  nor NOR2_642(G2868,G2798,G1232);
  nor NOR2_643(G2872,G2806,G2807);
  nor NOR2_644(G2875,G2811,G2812);
  nor NOR2_645(G2878,G2816,G2817);
  nor NOR2_646(G2881,G2821,G2822);
  nor NOR2_647(G2884,G2826,G2827);
  nor NOR2_648(G2887,G2831,G2832);
  nor NOR2_649(G2890,G2836,G2837);
  nor NOR2_650(G2893,G2841,G2842);
  nor NOR2_651(G2896,G2846,G2847);
  nor NOR2_652(G2899,G2851,G2852);
  nor NOR2_653(G2902,G2856,G2853);
  nor NOR2_654(G2906,G2789,G2859);
  nor NOR2_655(G2907,G2859,G2786);
  nor NOR2_656(G2908,G2863,G2864);
  nor NOR2_657(G2911,G2865,G1184);
  nor NOR2_658(G2915,G2798,G2868);
  nor NOR2_659(G2916,G2868,G1232);
  nor NOR2_660(G2917,G2685,G2868);
  nor NOR2_661(G2920,G2872,G2803);
  nor NOR2_662(G2924,G2875,G2808);
  nor NOR2_663(G2928,G2878,G2813);
  nor NOR2_664(G2932,G2881,G2818);
  nor NOR2_665(G2936,G2884,G2823);
  nor NOR2_666(G2940,G2887,G2828);
  nor NOR2_667(G2944,G2890,G2833);
  nor NOR2_668(G2948,G2893,G2838);
  nor NOR2_669(G2952,G2896,G2843);
  nor NOR2_670(G2956,G2899,G2848);
  nor NOR2_671(G2960,G2856,G2902);
  nor NOR2_672(G2961,G2902,G2853);
  nor NOR2_673(G2962,G2906,G2907);
  nor NOR2_674(G2965,G2908,G1136);
  nor NOR2_675(G2969,G2865,G2911);
  nor NOR2_676(G2970,G2911,G1184);
  nor NOR2_677(G2971,G2734,G2911);
  nor NOR2_678(G2974,G2915,G2916);
  nor NOR2_679(G2977,G1280,G2917);
  nor NOR2_680(G2981,G2872,G2920);
  nor NOR2_681(G2982,G2920,G2803);
  nor NOR2_682(G2983,G2875,G2924);
  nor NOR2_683(G2984,G2924,G2808);
  nor NOR2_684(G2985,G2878,G2928);
  nor NOR2_685(G2986,G2928,G2813);
  nor NOR2_686(G2987,G2881,G2932);
  nor NOR2_687(G2988,G2932,G2818);
  nor NOR2_688(G2989,G2884,G2936);
  nor NOR2_689(G2990,G2936,G2823);
  nor NOR2_690(G2991,G2887,G2940);
  nor NOR2_691(G2992,G2940,G2828);
  nor NOR2_692(G2993,G2890,G2944);
  nor NOR2_693(G2994,G2944,G2833);
  nor NOR2_694(G2995,G2893,G2948);
  nor NOR2_695(G2996,G2948,G2838);
  nor NOR2_696(G2997,G2896,G2952);
  nor NOR2_697(G2998,G2952,G2843);
  nor NOR2_698(G2999,G2899,G2956);
  nor NOR2_699(G3000,G2956,G2848);
  nor NOR2_700(G3001,G2960,G2961);
  nor NOR2_701(G3004,G2962,G1088);
  nor NOR2_702(G3008,G2908,G2965);
  nor NOR2_703(G3009,G2965,G1136);
  nor NOR2_704(G3010,G2792,G2965);
  nor NOR2_705(G3013,G2969,G2970);
  nor NOR2_706(G3016,G2974,G2971);
  nor NOR2_707(G3020,G1280,G2977);
  nor NOR2_708(G3021,G2977,G2917);
  nor NOR2_709(G3022,G2981,G2982);
  nor NOR2_710(G3025,G2983,G2984);
  nor NOR2_711(G3028,G2985,G2986);
  nor NOR2_712(G3031,G2987,G2988);
  nor NOR2_713(G3034,G2989,G2990);
  nor NOR2_714(G3037,G2991,G2992);
  nor NOR2_715(G3040,G2993,G2994);
  nor NOR2_716(G3043,G2995,G2996);
  nor NOR2_717(G3046,G2997,G2998);
  nor NOR2_718(G3049,G2999,G3000);
  nor NOR2_719(G3052,G3001,G1040);
  nor NOR2_720(G3056,G2962,G3004);
  nor NOR2_721(G3057,G3004,G1088);
  nor NOR2_722(G3058,G2859,G3004);
  nor NOR2_723(G3061,G3008,G3009);
  nor NOR2_724(G3064,G3013,G3010);
  nor NOR2_725(G3068,G2974,G3016);
  nor NOR2_726(G3069,G3016,G2971);
  nor NOR2_727(G3070,G3020,G3021);
  nor NOR2_728(G3073,G3022,G560);
  nor NOR2_729(G3077,G3025,G608);
  nor NOR2_730(G3081,G3028,G656);
  nor NOR2_731(G3085,G3031,G704);
  nor NOR2_732(G3089,G3034,G752);
  nor NOR2_733(G3093,G3037,G800);
  nor NOR2_734(G3097,G3040,G848);
  nor NOR2_735(G3101,G3043,G896);
  nor NOR2_736(G3105,G3046,G944);
  nor NOR2_737(G3109,G3049,G992);
  nor NOR2_738(G3113,G3001,G3052);
  nor NOR2_739(G3114,G3052,G1040);
  nor NOR2_740(G3115,G2902,G3052);
  nor NOR2_741(G3118,G3056,G3057);
  nor NOR2_742(G3121,G3061,G3058);
  nor NOR2_743(G3125,G3013,G3064);
  nor NOR2_744(G3126,G3064,G3010);
  nor NOR2_745(G3127,G3068,G3069);
  nor NOR2_746(G3130,G3070,G1235);
  nor NOR2_747(G3134,G3022,G3073);
  nor NOR2_748(G3135,G3073,G560);
  nor NOR2_749(G3136,G2920,G3073);
  nor NOR2_750(G3139,G3025,G3077);
  nor NOR2_751(G3140,G3077,G608);
  nor NOR2_752(G3141,G2924,G3077);
  nor NOR2_753(G3144,G3028,G3081);
  nor NOR2_754(G3145,G3081,G656);
  nor NOR2_755(G3146,G2928,G3081);
  nor NOR2_756(G3149,G3031,G3085);
  nor NOR2_757(G3150,G3085,G704);
  nor NOR2_758(G3151,G2932,G3085);
  nor NOR2_759(G3154,G3034,G3089);
  nor NOR2_760(G3155,G3089,G752);
  nor NOR2_761(G3156,G2936,G3089);
  nor NOR2_762(G3159,G3037,G3093);
  nor NOR2_763(G3160,G3093,G800);
  nor NOR2_764(G3161,G2940,G3093);
  nor NOR2_765(G3164,G3040,G3097);
  nor NOR2_766(G3165,G3097,G848);
  nor NOR2_767(G3166,G2944,G3097);
  nor NOR2_768(G3169,G3043,G3101);
  nor NOR2_769(G3170,G3101,G896);
  nor NOR2_770(G3171,G2948,G3101);
  nor NOR2_771(G3174,G3046,G3105);
  nor NOR2_772(G3175,G3105,G944);
  nor NOR2_773(G3176,G2952,G3105);
  nor NOR2_774(G3179,G3049,G3109);
  nor NOR2_775(G3180,G3109,G992);
  nor NOR2_776(G3181,G2956,G3109);
  nor NOR2_777(G3184,G3113,G3114);
  nor NOR2_778(G3187,G3118,G3115);
  nor NOR2_779(G3191,G3061,G3121);
  nor NOR2_780(G3192,G3121,G3058);
  nor NOR2_781(G3193,G3125,G3126);
  nor NOR2_782(G3196,G3127,G1187);
  nor NOR2_783(G3200,G3070,G3130);
  nor NOR2_784(G3201,G3130,G1235);
  nor NOR2_785(G3202,G2977,G3130);
  nor NOR2_786(G3205,G3139,G3140);
  nor NOR2_787(G3208,G3144,G3145);
  nor NOR2_788(G3211,G3149,G3150);
  nor NOR2_789(G3214,G3154,G3155);
  nor NOR2_790(G3217,G3159,G3160);
  nor NOR2_791(G3220,G3164,G3165);
  nor NOR2_792(G3223,G3169,G3170);
  nor NOR2_793(G3226,G3174,G3175);
  nor NOR2_794(G3229,G3179,G3180);
  nor NOR2_795(G3232,G3184,G3181);
  nor NOR2_796(G3236,G3118,G3187);
  nor NOR2_797(G3237,G3187,G3115);
  nor NOR2_798(G3238,G3191,G3192);
  nor NOR2_799(G3241,G3193,G1139);
  nor NOR2_800(G3245,G3127,G3196);
  nor NOR2_801(G3246,G3196,G1187);
  nor NOR2_802(G3247,G3016,G3196);
  nor NOR2_803(G3250,G3200,G3201);
  nor NOR2_804(G3253,G1283,G3202);
  nor NOR2_805(G3257,G3205,G3136);
  nor NOR2_806(G3261,G3208,G3141);
  nor NOR2_807(G3265,G3211,G3146);
  nor NOR2_808(G3269,G3214,G3151);
  nor NOR2_809(G3273,G3217,G3156);
  nor NOR2_810(G3277,G3220,G3161);
  nor NOR2_811(G3281,G3223,G3166);
  nor NOR2_812(G3285,G3226,G3171);
  nor NOR2_813(G3289,G3229,G3176);
  nor NOR2_814(G3293,G3184,G3232);
  nor NOR2_815(G3294,G3232,G3181);
  nor NOR2_816(G3295,G3236,G3237);
  nor NOR2_817(G3298,G3238,G1091);
  nor NOR2_818(G3302,G3193,G3241);
  nor NOR2_819(G3303,G3241,G1139);
  nor NOR2_820(G3304,G3064,G3241);
  nor NOR2_821(G3307,G3245,G3246);
  nor NOR2_822(G3310,G3250,G3247);
  nor NOR2_823(G3314,G1283,G3253);
  nor NOR2_824(G3315,G3253,G3202);
  nor NOR2_825(G3316,G3205,G3257);
  nor NOR2_826(G3317,G3257,G3136);
  nor NOR2_827(G3318,G3208,G3261);
  nor NOR2_828(G3319,G3261,G3141);
  nor NOR2_829(G3320,G3211,G3265);
  nor NOR2_830(G3321,G3265,G3146);
  nor NOR2_831(G3322,G3214,G3269);
  nor NOR2_832(G3323,G3269,G3151);
  nor NOR2_833(G3324,G3217,G3273);
  nor NOR2_834(G3325,G3273,G3156);
  nor NOR2_835(G3326,G3220,G3277);
  nor NOR2_836(G3327,G3277,G3161);
  nor NOR2_837(G3328,G3223,G3281);
  nor NOR2_838(G3329,G3281,G3166);
  nor NOR2_839(G3330,G3226,G3285);
  nor NOR2_840(G3331,G3285,G3171);
  nor NOR2_841(G3332,G3229,G3289);
  nor NOR2_842(G3333,G3289,G3176);
  nor NOR2_843(G3334,G3293,G3294);
  nor NOR2_844(G3337,G3295,G1043);
  nor NOR2_845(G3341,G3238,G3298);
  nor NOR2_846(G3342,G3298,G1091);
  nor NOR2_847(G3343,G3121,G3298);
  nor NOR2_848(G3346,G3302,G3303);
  nor NOR2_849(G3349,G3307,G3304);
  nor NOR2_850(G3353,G3250,G3310);
  nor NOR2_851(G3354,G3310,G3247);
  nor NOR2_852(G3355,G3314,G3315);
  nor NOR2_853(G3358,G3316,G3317);
  nor NOR2_854(G3361,G3318,G3319);
  nor NOR2_855(G3364,G3320,G3321);
  nor NOR2_856(G3367,G3322,G3323);
  nor NOR2_857(G3370,G3324,G3325);
  nor NOR2_858(G3373,G3326,G3327);
  nor NOR2_859(G3376,G3328,G3329);
  nor NOR2_860(G3379,G3330,G3331);
  nor NOR2_861(G3382,G3332,G3333);
  nor NOR2_862(G3385,G3334,G995);
  nor NOR2_863(G3389,G3295,G3337);
  nor NOR2_864(G3390,G3337,G1043);
  nor NOR2_865(G3391,G3187,G3337);
  nor NOR2_866(G3394,G3341,G3342);
  nor NOR2_867(G3397,G3346,G3343);
  nor NOR2_868(G3401,G3307,G3349);
  nor NOR2_869(G3402,G3349,G3304);
  nor NOR2_870(G3403,G3353,G3354);
  nor NOR2_871(G3406,G3355,G1238);
  nor NOR2_872(G3410,G3358,G563);
  nor NOR2_873(G3414,G3361,G611);
  nor NOR2_874(G3418,G3364,G659);
  nor NOR2_875(G3422,G3367,G707);
  nor NOR2_876(G3426,G3370,G755);
  nor NOR2_877(G3430,G3373,G803);
  nor NOR2_878(G3434,G3376,G851);
  nor NOR2_879(G3438,G3379,G899);
  nor NOR2_880(G3442,G3382,G947);
  nor NOR2_881(G3446,G3334,G3385);
  nor NOR2_882(G3447,G3385,G995);
  nor NOR2_883(G3448,G3232,G3385);
  nor NOR2_884(G3451,G3389,G3390);
  nor NOR2_885(G3454,G3394,G3391);
  nor NOR2_886(G3458,G3346,G3397);
  nor NOR2_887(G3459,G3397,G3343);
  nor NOR2_888(G3460,G3401,G3402);
  nor NOR2_889(G3463,G3403,G1190);
  nor NOR2_890(G3467,G3355,G3406);
  nor NOR2_891(G3468,G3406,G1238);
  nor NOR2_892(G3469,G3253,G3406);
  nor NOR2_893(G3472,G3358,G3410);
  nor NOR2_894(G3473,G3410,G563);
  nor NOR2_895(G3474,G3257,G3410);
  nor NOR2_896(G3477,G3361,G3414);
  nor NOR2_897(G3478,G3414,G611);
  nor NOR2_898(G3479,G3261,G3414);
  nor NOR2_899(G3482,G3364,G3418);
  nor NOR2_900(G3483,G3418,G659);
  nor NOR2_901(G3484,G3265,G3418);
  nor NOR2_902(G3487,G3367,G3422);
  nor NOR2_903(G3488,G3422,G707);
  nor NOR2_904(G3489,G3269,G3422);
  nor NOR2_905(G3492,G3370,G3426);
  nor NOR2_906(G3493,G3426,G755);
  nor NOR2_907(G3494,G3273,G3426);
  nor NOR2_908(G3497,G3373,G3430);
  nor NOR2_909(G3498,G3430,G803);
  nor NOR2_910(G3499,G3277,G3430);
  nor NOR2_911(G3502,G3376,G3434);
  nor NOR2_912(G3503,G3434,G851);
  nor NOR2_913(G3504,G3281,G3434);
  nor NOR2_914(G3507,G3379,G3438);
  nor NOR2_915(G3508,G3438,G899);
  nor NOR2_916(G3509,G3285,G3438);
  nor NOR2_917(G3512,G3382,G3442);
  nor NOR2_918(G3513,G3442,G947);
  nor NOR2_919(G3514,G3289,G3442);
  nor NOR2_920(G3517,G3446,G3447);
  nor NOR2_921(G3520,G3451,G3448);
  nor NOR2_922(G3524,G3394,G3454);
  nor NOR2_923(G3525,G3454,G3391);
  nor NOR2_924(G3526,G3458,G3459);
  nor NOR2_925(G3529,G3460,G1142);
  nor NOR2_926(G3533,G3403,G3463);
  nor NOR2_927(G3534,G3463,G1190);
  nor NOR2_928(G3535,G3310,G3463);
  nor NOR2_929(G3538,G3467,G3468);
  nor NOR2_930(G3541,G1286,G3469);
  nor NOR2_931(G3545,G3477,G3478);
  nor NOR2_932(G3548,G3482,G3483);
  nor NOR2_933(G3551,G3487,G3488);
  nor NOR2_934(G3554,G3492,G3493);
  nor NOR2_935(G3557,G3497,G3498);
  nor NOR2_936(G3560,G3502,G3503);
  nor NOR2_937(G3563,G3507,G3508);
  nor NOR2_938(G3566,G3512,G3513);
  nor NOR2_939(G3569,G3517,G3514);
  nor NOR2_940(G3573,G3451,G3520);
  nor NOR2_941(G3574,G3520,G3448);
  nor NOR2_942(G3575,G3524,G3525);
  nor NOR2_943(G3578,G3526,G1094);
  nor NOR2_944(G3582,G3460,G3529);
  nor NOR2_945(G3583,G3529,G1142);
  nor NOR2_946(G3584,G3349,G3529);
  nor NOR2_947(G3587,G3533,G3534);
  nor NOR2_948(G3590,G3538,G3535);
  nor NOR2_949(G3594,G1286,G3541);
  nor NOR2_950(G3595,G3541,G3469);
  nor NOR2_951(G3596,G3545,G3474);
  nor NOR2_952(G3600,G3548,G3479);
  nor NOR2_953(G3604,G3551,G3484);
  nor NOR2_954(G3608,G3554,G3489);
  nor NOR2_955(G3612,G3557,G3494);
  nor NOR2_956(G3616,G3560,G3499);
  nor NOR2_957(G3620,G3563,G3504);
  nor NOR2_958(G3624,G3566,G3509);
  nor NOR2_959(G3628,G3517,G3569);
  nor NOR2_960(G3629,G3569,G3514);
  nor NOR2_961(G3630,G3573,G3574);
  nor NOR2_962(G3633,G3575,G1046);
  nor NOR2_963(G3637,G3526,G3578);
  nor NOR2_964(G3638,G3578,G1094);
  nor NOR2_965(G3639,G3397,G3578);
  nor NOR2_966(G3642,G3582,G3583);
  nor NOR2_967(G3645,G3587,G3584);
  nor NOR2_968(G3649,G3538,G3590);
  nor NOR2_969(G3650,G3590,G3535);
  nor NOR2_970(G3651,G3594,G3595);
  nor NOR2_971(G3654,G3545,G3596);
  nor NOR2_972(G3655,G3596,G3474);
  nor NOR2_973(G3656,G3548,G3600);
  nor NOR2_974(G3657,G3600,G3479);
  nor NOR2_975(G3658,G3551,G3604);
  nor NOR2_976(G3659,G3604,G3484);
  nor NOR2_977(G3660,G3554,G3608);
  nor NOR2_978(G3661,G3608,G3489);
  nor NOR2_979(G3662,G3557,G3612);
  nor NOR2_980(G3663,G3612,G3494);
  nor NOR2_981(G3664,G3560,G3616);
  nor NOR2_982(G3665,G3616,G3499);
  nor NOR2_983(G3666,G3563,G3620);
  nor NOR2_984(G3667,G3620,G3504);
  nor NOR2_985(G3668,G3566,G3624);
  nor NOR2_986(G3669,G3624,G3509);
  nor NOR2_987(G3670,G3628,G3629);
  nor NOR2_988(G3673,G3630,G998);
  nor NOR2_989(G3677,G3575,G3633);
  nor NOR2_990(G3678,G3633,G1046);
  nor NOR2_991(G3679,G3454,G3633);
  nor NOR2_992(G3682,G3637,G3638);
  nor NOR2_993(G3685,G3642,G3639);
  nor NOR2_994(G3689,G3587,G3645);
  nor NOR2_995(G3690,G3645,G3584);
  nor NOR2_996(G3691,G3649,G3650);
  nor NOR2_997(G3694,G3651,G1241);
  nor NOR2_998(G3698,G3654,G3655);
  nor NOR2_999(G3701,G3656,G3657);
  nor NOR2_1000(G3704,G3658,G3659);
  nor NOR2_1001(G3707,G3660,G3661);
  nor NOR2_1002(G3710,G3662,G3663);
  nor NOR2_1003(G3713,G3664,G3665);
  nor NOR2_1004(G3716,G3666,G3667);
  nor NOR2_1005(G3719,G3668,G3669);
  nor NOR2_1006(G3722,G3670,G950);
  nor NOR2_1007(G3726,G3630,G3673);
  nor NOR2_1008(G3727,G3673,G998);
  nor NOR2_1009(G3728,G3520,G3673);
  nor NOR2_1010(G3731,G3677,G3678);
  nor NOR2_1011(G3734,G3682,G3679);
  nor NOR2_1012(G3738,G3642,G3685);
  nor NOR2_1013(G3739,G3685,G3639);
  nor NOR2_1014(G3740,G3689,G3690);
  nor NOR2_1015(G3743,G3691,G1193);
  nor NOR2_1016(G3747,G3651,G3694);
  nor NOR2_1017(G3748,G3694,G1241);
  nor NOR2_1018(G3749,G3541,G3694);
  nor NOR2_1019(G3752,G3698,G566);
  nor NOR2_1020(G3756,G3701,G614);
  nor NOR2_1021(G3760,G3704,G662);
  nor NOR2_1022(G3764,G3707,G710);
  nor NOR2_1023(G3768,G3710,G758);
  nor NOR2_1024(G3772,G3713,G806);
  nor NOR2_1025(G3776,G3716,G854);
  nor NOR2_1026(G3780,G3719,G902);
  nor NOR2_1027(G3784,G3670,G3722);
  nor NOR2_1028(G3785,G3722,G950);
  nor NOR2_1029(G3786,G3569,G3722);
  nor NOR2_1030(G3789,G3726,G3727);
  nor NOR2_1031(G3792,G3731,G3728);
  nor NOR2_1032(G3796,G3682,G3734);
  nor NOR2_1033(G3797,G3734,G3679);
  nor NOR2_1034(G3798,G3738,G3739);
  nor NOR2_1035(G3801,G3740,G1145);
  nor NOR2_1036(G3805,G3691,G3743);
  nor NOR2_1037(G3806,G3743,G1193);
  nor NOR2_1038(G3807,G3590,G3743);
  nor NOR2_1039(G3810,G3747,G3748);
  nor NOR2_1040(G3813,G1289,G3749);
  nor NOR2_1041(G3817,G3698,G3752);
  nor NOR2_1042(G3818,G3752,G566);
  nor NOR2_1043(G3819,G3596,G3752);
  nor NOR2_1044(G3822,G3701,G3756);
  nor NOR2_1045(G3823,G3756,G614);
  nor NOR2_1046(G3824,G3600,G3756);
  nor NOR2_1047(G3827,G3704,G3760);
  nor NOR2_1048(G3828,G3760,G662);
  nor NOR2_1049(G3829,G3604,G3760);
  nor NOR2_1050(G3832,G3707,G3764);
  nor NOR2_1051(G3833,G3764,G710);
  nor NOR2_1052(G3834,G3608,G3764);
  nor NOR2_1053(G3837,G3710,G3768);
  nor NOR2_1054(G3838,G3768,G758);
  nor NOR2_1055(G3839,G3612,G3768);
  nor NOR2_1056(G3842,G3713,G3772);
  nor NOR2_1057(G3843,G3772,G806);
  nor NOR2_1058(G3844,G3616,G3772);
  nor NOR2_1059(G3847,G3716,G3776);
  nor NOR2_1060(G3848,G3776,G854);
  nor NOR2_1061(G3849,G3620,G3776);
  nor NOR2_1062(G3852,G3719,G3780);
  nor NOR2_1063(G3853,G3780,G902);
  nor NOR2_1064(G3854,G3624,G3780);
  nor NOR2_1065(G3857,G3784,G3785);
  nor NOR2_1066(G3860,G3789,G3786);
  nor NOR2_1067(G3864,G3731,G3792);
  nor NOR2_1068(G3865,G3792,G3728);
  nor NOR2_1069(G3866,G3796,G3797);
  nor NOR2_1070(G3869,G3798,G1097);
  nor NOR2_1071(G3873,G3740,G3801);
  nor NOR2_1072(G3874,G3801,G1145);
  nor NOR2_1073(G3875,G3645,G3801);
  nor NOR2_1074(G3878,G3805,G3806);
  nor NOR2_1075(G3881,G3810,G3807);
  nor NOR2_1076(G3885,G1289,G3813);
  nor NOR2_1077(G3886,G3813,G3749);
  nor NOR2_1078(G3887,G3822,G3823);
  nor NOR2_1079(G3890,G3827,G3828);
  nor NOR2_1080(G3893,G3832,G3833);
  nor NOR2_1081(G3896,G3837,G3838);
  nor NOR2_1082(G3899,G3842,G3843);
  nor NOR2_1083(G3902,G3847,G3848);
  nor NOR2_1084(G3905,G3852,G3853);
  nor NOR2_1085(G3908,G3857,G3854);
  nor NOR2_1086(G3912,G3789,G3860);
  nor NOR2_1087(G3913,G3860,G3786);
  nor NOR2_1088(G3914,G3864,G3865);
  nor NOR2_1089(G3917,G3866,G1049);
  nor NOR2_1090(G3921,G3798,G3869);
  nor NOR2_1091(G3922,G3869,G1097);
  nor NOR2_1092(G3923,G3685,G3869);
  nor NOR2_1093(G3926,G3873,G3874);
  nor NOR2_1094(G3929,G3878,G3875);
  nor NOR2_1095(G3933,G3810,G3881);
  nor NOR2_1096(G3934,G3881,G3807);
  nor NOR2_1097(G3935,G3885,G3886);
  nor NOR2_1098(G3938,G3887,G3819);
  nor NOR2_1099(G3942,G3890,G3824);
  nor NOR2_1100(G3946,G3893,G3829);
  nor NOR2_1101(G3950,G3896,G3834);
  nor NOR2_1102(G3954,G3899,G3839);
  nor NOR2_1103(G3958,G3902,G3844);
  nor NOR2_1104(G3962,G3905,G3849);
  nor NOR2_1105(G3966,G3857,G3908);
  nor NOR2_1106(G3967,G3908,G3854);
  nor NOR2_1107(G3968,G3912,G3913);
  nor NOR2_1108(G3971,G3914,G1001);
  nor NOR2_1109(G3975,G3866,G3917);
  nor NOR2_1110(G3976,G3917,G1049);
  nor NOR2_1111(G3977,G3734,G3917);
  nor NOR2_1112(G3980,G3921,G3922);
  nor NOR2_1113(G3983,G3926,G3923);
  nor NOR2_1114(G3987,G3878,G3929);
  nor NOR2_1115(G3988,G3929,G3875);
  nor NOR2_1116(G3989,G3933,G3934);
  nor NOR2_1117(G3992,G3935,G1244);
  nor NOR2_1118(G3996,G3887,G3938);
  nor NOR2_1119(G3997,G3938,G3819);
  nor NOR2_1120(G3998,G3890,G3942);
  nor NOR2_1121(G3999,G3942,G3824);
  nor NOR2_1122(G4000,G3893,G3946);
  nor NOR2_1123(G4001,G3946,G3829);
  nor NOR2_1124(G4002,G3896,G3950);
  nor NOR2_1125(G4003,G3950,G3834);
  nor NOR2_1126(G4004,G3899,G3954);
  nor NOR2_1127(G4005,G3954,G3839);
  nor NOR2_1128(G4006,G3902,G3958);
  nor NOR2_1129(G4007,G3958,G3844);
  nor NOR2_1130(G4008,G3905,G3962);
  nor NOR2_1131(G4009,G3962,G3849);
  nor NOR2_1132(G4010,G3966,G3967);
  nor NOR2_1133(G4013,G3968,G953);
  nor NOR2_1134(G4017,G3914,G3971);
  nor NOR2_1135(G4018,G3971,G1001);
  nor NOR2_1136(G4019,G3792,G3971);
  nor NOR2_1137(G4022,G3975,G3976);
  nor NOR2_1138(G4025,G3980,G3977);
  nor NOR2_1139(G4029,G3926,G3983);
  nor NOR2_1140(G4030,G3983,G3923);
  nor NOR2_1141(G4031,G3987,G3988);
  nor NOR2_1142(G4034,G3989,G1196);
  nor NOR2_1143(G4038,G3935,G3992);
  nor NOR2_1144(G4039,G3992,G1244);
  nor NOR2_1145(G4040,G3813,G3992);
  nor NOR2_1146(G4043,G3996,G3997);
  nor NOR2_1147(G4046,G3998,G3999);
  nor NOR2_1148(G4049,G4000,G4001);
  nor NOR2_1149(G4052,G4002,G4003);
  nor NOR2_1150(G4055,G4004,G4005);
  nor NOR2_1151(G4058,G4006,G4007);
  nor NOR2_1152(G4061,G4008,G4009);
  nor NOR2_1153(G4064,G4010,G905);
  nor NOR2_1154(G4068,G3968,G4013);
  nor NOR2_1155(G4069,G4013,G953);
  nor NOR2_1156(G4070,G3860,G4013);
  nor NOR2_1157(G4073,G4017,G4018);
  nor NOR2_1158(G4076,G4022,G4019);
  nor NOR2_1159(G4080,G3980,G4025);
  nor NOR2_1160(G4081,G4025,G3977);
  nor NOR2_1161(G4082,G4029,G4030);
  nor NOR2_1162(G4085,G4031,G1148);
  nor NOR2_1163(G4089,G3989,G4034);
  nor NOR2_1164(G4090,G4034,G1196);
  nor NOR2_1165(G4091,G3881,G4034);
  nor NOR2_1166(G4094,G4038,G4039);
  nor NOR2_1167(G4097,G1292,G4040);
  nor NOR2_1168(G4101,G4043,G569);
  nor NOR2_1169(G4105,G4046,G617);
  nor NOR2_1170(G4109,G4049,G665);
  nor NOR2_1171(G4113,G4052,G713);
  nor NOR2_1172(G4117,G4055,G761);
  nor NOR2_1173(G4121,G4058,G809);
  nor NOR2_1174(G4125,G4061,G857);
  nor NOR2_1175(G4129,G4010,G4064);
  nor NOR2_1176(G4130,G4064,G905);
  nor NOR2_1177(G4131,G3908,G4064);
  nor NOR2_1178(G4134,G4068,G4069);
  nor NOR2_1179(G4137,G4073,G4070);
  nor NOR2_1180(G4141,G4022,G4076);
  nor NOR2_1181(G4142,G4076,G4019);
  nor NOR2_1182(G4143,G4080,G4081);
  nor NOR2_1183(G4146,G4082,G1100);
  nor NOR2_1184(G4150,G4031,G4085);
  nor NOR2_1185(G4151,G4085,G1148);
  nor NOR2_1186(G4152,G3929,G4085);
  nor NOR2_1187(G4155,G4089,G4090);
  nor NOR2_1188(G4158,G4094,G4091);
  nor NOR2_1189(G4162,G1292,G4097);
  nor NOR2_1190(G4163,G4097,G4040);
  nor NOR2_1191(G4164,G4043,G4101);
  nor NOR2_1192(G4165,G4101,G569);
  nor NOR2_1193(G4166,G3938,G4101);
  nor NOR2_1194(G4169,G4046,G4105);
  nor NOR2_1195(G4170,G4105,G617);
  nor NOR2_1196(G4171,G3942,G4105);
  nor NOR2_1197(G4174,G4049,G4109);
  nor NOR2_1198(G4175,G4109,G665);
  nor NOR2_1199(G4176,G3946,G4109);
  nor NOR2_1200(G4179,G4052,G4113);
  nor NOR2_1201(G4180,G4113,G713);
  nor NOR2_1202(G4181,G3950,G4113);
  nor NOR2_1203(G4184,G4055,G4117);
  nor NOR2_1204(G4185,G4117,G761);
  nor NOR2_1205(G4186,G3954,G4117);
  nor NOR2_1206(G4189,G4058,G4121);
  nor NOR2_1207(G4190,G4121,G809);
  nor NOR2_1208(G4191,G3958,G4121);
  nor NOR2_1209(G4194,G4061,G4125);
  nor NOR2_1210(G4195,G4125,G857);
  nor NOR2_1211(G4196,G3962,G4125);
  nor NOR2_1212(G4199,G4129,G4130);
  nor NOR2_1213(G4202,G4134,G4131);
  nor NOR2_1214(G4206,G4073,G4137);
  nor NOR2_1215(G4207,G4137,G4070);
  nor NOR2_1216(G4208,G4141,G4142);
  nor NOR2_1217(G4211,G4143,G1052);
  nor NOR2_1218(G4215,G4082,G4146);
  nor NOR2_1219(G4216,G4146,G1100);
  nor NOR2_1220(G4217,G3983,G4146);
  nor NOR2_1221(G4220,G4150,G4151);
  nor NOR2_1222(G4223,G4155,G4152);
  nor NOR2_1223(G4227,G4094,G4158);
  nor NOR2_1224(G4228,G4158,G4091);
  nor NOR2_1225(G4229,G4162,G4163);
  nor NOR2_1226(G4232,G4169,G4170);
  nor NOR2_1227(G4235,G4174,G4175);
  nor NOR2_1228(G4238,G4179,G4180);
  nor NOR2_1229(G4241,G4184,G4185);
  nor NOR2_1230(G4244,G4189,G4190);
  nor NOR2_1231(G4247,G4194,G4195);
  nor NOR2_1232(G4250,G4199,G4196);
  nor NOR2_1233(G4254,G4134,G4202);
  nor NOR2_1234(G4255,G4202,G4131);
  nor NOR2_1235(G4256,G4206,G4207);
  nor NOR2_1236(G4259,G4208,G1004);
  nor NOR2_1237(G4263,G4143,G4211);
  nor NOR2_1238(G4264,G4211,G1052);
  nor NOR2_1239(G4265,G4025,G4211);
  nor NOR2_1240(G4268,G4215,G4216);
  nor NOR2_1241(G4271,G4220,G4217);
  nor NOR2_1242(G4275,G4155,G4223);
  nor NOR2_1243(G4276,G4223,G4152);
  nor NOR2_1244(G4277,G4227,G4228);
  nor NOR2_1245(G4280,G4229,G1247);
  nor NOR2_1246(G4284,G4232,G4166);
  nor NOR2_1247(G4288,G4235,G4171);
  nor NOR2_1248(G4292,G4238,G4176);
  nor NOR2_1249(G4296,G4241,G4181);
  nor NOR2_1250(G4300,G4244,G4186);
  nor NOR2_1251(G4304,G4247,G4191);
  nor NOR2_1252(G4308,G4199,G4250);
  nor NOR2_1253(G4309,G4250,G4196);
  nor NOR2_1254(G4310,G4254,G4255);
  nor NOR2_1255(G4313,G4256,G956);
  nor NOR2_1256(G4317,G4208,G4259);
  nor NOR2_1257(G4318,G4259,G1004);
  nor NOR2_1258(G4319,G4076,G4259);
  nor NOR2_1259(G4322,G4263,G4264);
  nor NOR2_1260(G4325,G4268,G4265);
  nor NOR2_1261(G4329,G4220,G4271);
  nor NOR2_1262(G4330,G4271,G4217);
  nor NOR2_1263(G4331,G4275,G4276);
  nor NOR2_1264(G4334,G4277,G1199);
  nor NOR2_1265(G4338,G4229,G4280);
  nor NOR2_1266(G4339,G4280,G1247);
  nor NOR2_1267(G4340,G4097,G4280);
  nor NOR2_1268(G4343,G4232,G4284);
  nor NOR2_1269(G4344,G4284,G4166);
  nor NOR2_1270(G4345,G4235,G4288);
  nor NOR2_1271(G4346,G4288,G4171);
  nor NOR2_1272(G4347,G4238,G4292);
  nor NOR2_1273(G4348,G4292,G4176);
  nor NOR2_1274(G4349,G4241,G4296);
  nor NOR2_1275(G4350,G4296,G4181);
  nor NOR2_1276(G4351,G4244,G4300);
  nor NOR2_1277(G4352,G4300,G4186);
  nor NOR2_1278(G4353,G4247,G4304);
  nor NOR2_1279(G4354,G4304,G4191);
  nor NOR2_1280(G4355,G4308,G4309);
  nor NOR2_1281(G4358,G4310,G908);
  nor NOR2_1282(G4362,G4256,G4313);
  nor NOR2_1283(G4363,G4313,G956);
  nor NOR2_1284(G4364,G4137,G4313);
  nor NOR2_1285(G4367,G4317,G4318);
  nor NOR2_1286(G4370,G4322,G4319);
  nor NOR2_1287(G4374,G4268,G4325);
  nor NOR2_1288(G4375,G4325,G4265);
  nor NOR2_1289(G4376,G4329,G4330);
  nor NOR2_1290(G4379,G4331,G1151);
  nor NOR2_1291(G4383,G4277,G4334);
  nor NOR2_1292(G4384,G4334,G1199);
  nor NOR2_1293(G4385,G4158,G4334);
  nor NOR2_1294(G4388,G4338,G4339);
  nor NOR2_1295(G4391,G1295,G4340);
  nor NOR2_1296(G4395,G4343,G4344);
  nor NOR2_1297(G4398,G4345,G4346);
  nor NOR2_1298(G4401,G4347,G4348);
  nor NOR2_1299(G4404,G4349,G4350);
  nor NOR2_1300(G4407,G4351,G4352);
  nor NOR2_1301(G4410,G4353,G4354);
  nor NOR2_1302(G4413,G4355,G860);
  nor NOR2_1303(G4417,G4310,G4358);
  nor NOR2_1304(G4418,G4358,G908);
  nor NOR2_1305(G4419,G4202,G4358);
  nor NOR2_1306(G4422,G4362,G4363);
  nor NOR2_1307(G4425,G4367,G4364);
  nor NOR2_1308(G4429,G4322,G4370);
  nor NOR2_1309(G4430,G4370,G4319);
  nor NOR2_1310(G4431,G4374,G4375);
  nor NOR2_1311(G4434,G4376,G1103);
  nor NOR2_1312(G4438,G4331,G4379);
  nor NOR2_1313(G4439,G4379,G1151);
  nor NOR2_1314(G4440,G4223,G4379);
  nor NOR2_1315(G4443,G4383,G4384);
  nor NOR2_1316(G4446,G4388,G4385);
  nor NOR2_1317(G4450,G1295,G4391);
  nor NOR2_1318(G4451,G4391,G4340);
  nor NOR2_1319(G4452,G4395,G572);
  nor NOR2_1320(G4456,G4398,G620);
  nor NOR2_1321(G4460,G4401,G668);
  nor NOR2_1322(G4464,G4404,G716);
  nor NOR2_1323(G4468,G4407,G764);
  nor NOR2_1324(G4472,G4410,G812);
  nor NOR2_1325(G4476,G4355,G4413);
  nor NOR2_1326(G4477,G4413,G860);
  nor NOR2_1327(G4478,G4250,G4413);
  nor NOR2_1328(G4481,G4417,G4418);
  nor NOR2_1329(G4484,G4422,G4419);
  nor NOR2_1330(G4488,G4367,G4425);
  nor NOR2_1331(G4489,G4425,G4364);
  nor NOR2_1332(G4490,G4429,G4430);
  nor NOR2_1333(G4493,G4431,G1055);
  nor NOR2_1334(G4497,G4376,G4434);
  nor NOR2_1335(G4498,G4434,G1103);
  nor NOR2_1336(G4499,G4271,G4434);
  nor NOR2_1337(G4502,G4438,G4439);
  nor NOR2_1338(G4505,G4443,G4440);
  nor NOR2_1339(G4509,G4388,G4446);
  nor NOR2_1340(G4510,G4446,G4385);
  nor NOR2_1341(G4511,G4450,G4451);
  nor NOR2_1342(G4514,G4395,G4452);
  nor NOR2_1343(G4515,G4452,G572);
  nor NOR2_1344(G4516,G4284,G4452);
  nor NOR2_1345(G4519,G4398,G4456);
  nor NOR2_1346(G4520,G4456,G620);
  nor NOR2_1347(G4521,G4288,G4456);
  nor NOR2_1348(G4524,G4401,G4460);
  nor NOR2_1349(G4525,G4460,G668);
  nor NOR2_1350(G4526,G4292,G4460);
  nor NOR2_1351(G4529,G4404,G4464);
  nor NOR2_1352(G4530,G4464,G716);
  nor NOR2_1353(G4531,G4296,G4464);
  nor NOR2_1354(G4534,G4407,G4468);
  nor NOR2_1355(G4535,G4468,G764);
  nor NOR2_1356(G4536,G4300,G4468);
  nor NOR2_1357(G4539,G4410,G4472);
  nor NOR2_1358(G4540,G4472,G812);
  nor NOR2_1359(G4541,G4304,G4472);
  nor NOR2_1360(G4544,G4476,G4477);
  nor NOR2_1361(G4547,G4481,G4478);
  nor NOR2_1362(G4551,G4422,G4484);
  nor NOR2_1363(G4552,G4484,G4419);
  nor NOR2_1364(G4553,G4488,G4489);
  nor NOR2_1365(G4556,G4490,G1007);
  nor NOR2_1366(G4560,G4431,G4493);
  nor NOR2_1367(G4561,G4493,G1055);
  nor NOR2_1368(G4562,G4325,G4493);
  nor NOR2_1369(G4565,G4497,G4498);
  nor NOR2_1370(G4568,G4502,G4499);
  nor NOR2_1371(G4572,G4443,G4505);
  nor NOR2_1372(G4573,G4505,G4440);
  nor NOR2_1373(G4574,G4509,G4510);
  nor NOR2_1374(G4577,G4511,G1250);
  nor NOR2_1375(G4581,G4519,G4520);
  nor NOR2_1376(G4584,G4524,G4525);
  nor NOR2_1377(G4587,G4529,G4530);
  nor NOR2_1378(G4590,G4534,G4535);
  nor NOR2_1379(G4593,G4539,G4540);
  nor NOR2_1380(G4596,G4544,G4541);
  nor NOR2_1381(G4600,G4481,G4547);
  nor NOR2_1382(G4601,G4547,G4478);
  nor NOR2_1383(G4602,G4551,G4552);
  nor NOR2_1384(G4605,G4553,G959);
  nor NOR2_1385(G4609,G4490,G4556);
  nor NOR2_1386(G4610,G4556,G1007);
  nor NOR2_1387(G4611,G4370,G4556);
  nor NOR2_1388(G4614,G4560,G4561);
  nor NOR2_1389(G4617,G4565,G4562);
  nor NOR2_1390(G4621,G4502,G4568);
  nor NOR2_1391(G4622,G4568,G4499);
  nor NOR2_1392(G4623,G4572,G4573);
  nor NOR2_1393(G4626,G4574,G1202);
  nor NOR2_1394(G4630,G4511,G4577);
  nor NOR2_1395(G4631,G4577,G1250);
  nor NOR2_1396(G4632,G4391,G4577);
  nor NOR2_1397(G4635,G4581,G4516);
  nor NOR2_1398(G4639,G4584,G4521);
  nor NOR2_1399(G4643,G4587,G4526);
  nor NOR2_1400(G4647,G4590,G4531);
  nor NOR2_1401(G4651,G4593,G4536);
  nor NOR2_1402(G4655,G4544,G4596);
  nor NOR2_1403(G4656,G4596,G4541);
  nor NOR2_1404(G4657,G4600,G4601);
  nor NOR2_1405(G4660,G4602,G911);
  nor NOR2_1406(G4664,G4553,G4605);
  nor NOR2_1407(G4665,G4605,G959);
  nor NOR2_1408(G4666,G4425,G4605);
  nor NOR2_1409(G4669,G4609,G4610);
  nor NOR2_1410(G4672,G4614,G4611);
  nor NOR2_1411(G4676,G4565,G4617);
  nor NOR2_1412(G4677,G4617,G4562);
  nor NOR2_1413(G4678,G4621,G4622);
  nor NOR2_1414(G4681,G4623,G1154);
  nor NOR2_1415(G4685,G4574,G4626);
  nor NOR2_1416(G4686,G4626,G1202);
  nor NOR2_1417(G4687,G4446,G4626);
  nor NOR2_1418(G4690,G4630,G4631);
  nor NOR2_1419(G4693,G1298,G4632);
  nor NOR2_1420(G4697,G4581,G4635);
  nor NOR2_1421(G4698,G4635,G4516);
  nor NOR2_1422(G4699,G4584,G4639);
  nor NOR2_1423(G4700,G4639,G4521);
  nor NOR2_1424(G4701,G4587,G4643);
  nor NOR2_1425(G4702,G4643,G4526);
  nor NOR2_1426(G4703,G4590,G4647);
  nor NOR2_1427(G4704,G4647,G4531);
  nor NOR2_1428(G4705,G4593,G4651);
  nor NOR2_1429(G4706,G4651,G4536);
  nor NOR2_1430(G4707,G4655,G4656);
  nor NOR2_1431(G4710,G4657,G863);
  nor NOR2_1432(G4714,G4602,G4660);
  nor NOR2_1433(G4715,G4660,G911);
  nor NOR2_1434(G4716,G4484,G4660);
  nor NOR2_1435(G4719,G4664,G4665);
  nor NOR2_1436(G4722,G4669,G4666);
  nor NOR2_1437(G4726,G4614,G4672);
  nor NOR2_1438(G4727,G4672,G4611);
  nor NOR2_1439(G4728,G4676,G4677);
  nor NOR2_1440(G4731,G4678,G1106);
  nor NOR2_1441(G4735,G4623,G4681);
  nor NOR2_1442(G4736,G4681,G1154);
  nor NOR2_1443(G4737,G4505,G4681);
  nor NOR2_1444(G4740,G4685,G4686);
  nor NOR2_1445(G4743,G4690,G4687);
  nor NOR2_1446(G4747,G1298,G4693);
  nor NOR2_1447(G4748,G4693,G4632);
  nor NOR2_1448(G4749,G4697,G4698);
  nor NOR2_1449(G4752,G4699,G4700);
  nor NOR2_1450(G4755,G4701,G4702);
  nor NOR2_1451(G4758,G4703,G4704);
  nor NOR2_1452(G4761,G4705,G4706);
  nor NOR2_1453(G4764,G4707,G815);
  nor NOR2_1454(G4768,G4657,G4710);
  nor NOR2_1455(G4769,G4710,G863);
  nor NOR2_1456(G4770,G4547,G4710);
  nor NOR2_1457(G4773,G4714,G4715);
  nor NOR2_1458(G4776,G4719,G4716);
  nor NOR2_1459(G4780,G4669,G4722);
  nor NOR2_1460(G4781,G4722,G4666);
  nor NOR2_1461(G4782,G4726,G4727);
  nor NOR2_1462(G4785,G4728,G1058);
  nor NOR2_1463(G4789,G4678,G4731);
  nor NOR2_1464(G4790,G4731,G1106);
  nor NOR2_1465(G4791,G4568,G4731);
  nor NOR2_1466(G4794,G4735,G4736);
  nor NOR2_1467(G4797,G4740,G4737);
  nor NOR2_1468(G4801,G4690,G4743);
  nor NOR2_1469(G4802,G4743,G4687);
  nor NOR2_1470(G4803,G4747,G4748);
  nor NOR2_1471(G4806,G4749,G575);
  nor NOR2_1472(G4810,G4752,G623);
  nor NOR2_1473(G4814,G4755,G671);
  nor NOR2_1474(G4818,G4758,G719);
  nor NOR2_1475(G4822,G4761,G767);
  nor NOR2_1476(G4826,G4707,G4764);
  nor NOR2_1477(G4827,G4764,G815);
  nor NOR2_1478(G4828,G4596,G4764);
  nor NOR2_1479(G4831,G4768,G4769);
  nor NOR2_1480(G4834,G4773,G4770);
  nor NOR2_1481(G4838,G4719,G4776);
  nor NOR2_1482(G4839,G4776,G4716);
  nor NOR2_1483(G4840,G4780,G4781);
  nor NOR2_1484(G4843,G4782,G1010);
  nor NOR2_1485(G4847,G4728,G4785);
  nor NOR2_1486(G4848,G4785,G1058);
  nor NOR2_1487(G4849,G4617,G4785);
  nor NOR2_1488(G4852,G4789,G4790);
  nor NOR2_1489(G4855,G4794,G4791);
  nor NOR2_1490(G4859,G4740,G4797);
  nor NOR2_1491(G4860,G4797,G4737);
  nor NOR2_1492(G4861,G4801,G4802);
  nor NOR2_1493(G4864,G4803,G1253);
  nor NOR2_1494(G4868,G4749,G4806);
  nor NOR2_1495(G4869,G4806,G575);
  nor NOR2_1496(G4870,G4635,G4806);
  nor NOR2_1497(G4873,G4752,G4810);
  nor NOR2_1498(G4874,G4810,G623);
  nor NOR2_1499(G4875,G4639,G4810);
  nor NOR2_1500(G4878,G4755,G4814);
  nor NOR2_1501(G4879,G4814,G671);
  nor NOR2_1502(G4880,G4643,G4814);
  nor NOR2_1503(G4883,G4758,G4818);
  nor NOR2_1504(G4884,G4818,G719);
  nor NOR2_1505(G4885,G4647,G4818);
  nor NOR2_1506(G4888,G4761,G4822);
  nor NOR2_1507(G4889,G4822,G767);
  nor NOR2_1508(G4890,G4651,G4822);
  nor NOR2_1509(G4893,G4826,G4827);
  nor NOR2_1510(G4896,G4831,G4828);
  nor NOR2_1511(G4900,G4773,G4834);
  nor NOR2_1512(G4901,G4834,G4770);
  nor NOR2_1513(G4902,G4838,G4839);
  nor NOR2_1514(G4905,G4840,G962);
  nor NOR2_1515(G4909,G4782,G4843);
  nor NOR2_1516(G4910,G4843,G1010);
  nor NOR2_1517(G4911,G4672,G4843);
  nor NOR2_1518(G4914,G4847,G4848);
  nor NOR2_1519(G4917,G4852,G4849);
  nor NOR2_1520(G4921,G4794,G4855);
  nor NOR2_1521(G4922,G4855,G4791);
  nor NOR2_1522(G4923,G4859,G4860);
  nor NOR2_1523(G4926,G4861,G1205);
  nor NOR2_1524(G4930,G4803,G4864);
  nor NOR2_1525(G4931,G4864,G1253);
  nor NOR2_1526(G4932,G4693,G4864);
  nor NOR2_1527(G4935,G4873,G4874);
  nor NOR2_1528(G4938,G4878,G4879);
  nor NOR2_1529(G4941,G4883,G4884);
  nor NOR2_1530(G4944,G4888,G4889);
  nor NOR2_1531(G4947,G4893,G4890);
  nor NOR2_1532(G4951,G4831,G4896);
  nor NOR2_1533(G4952,G4896,G4828);
  nor NOR2_1534(G4953,G4900,G4901);
  nor NOR2_1535(G4956,G4902,G914);
  nor NOR2_1536(G4960,G4840,G4905);
  nor NOR2_1537(G4961,G4905,G962);
  nor NOR2_1538(G4962,G4722,G4905);
  nor NOR2_1539(G4965,G4909,G4910);
  nor NOR2_1540(G4968,G4914,G4911);
  nor NOR2_1541(G4972,G4852,G4917);
  nor NOR2_1542(G4973,G4917,G4849);
  nor NOR2_1543(G4974,G4921,G4922);
  nor NOR2_1544(G4977,G4923,G1157);
  nor NOR2_1545(G4981,G4861,G4926);
  nor NOR2_1546(G4982,G4926,G1205);
  nor NOR2_1547(G4983,G4743,G4926);
  nor NOR2_1548(G4986,G4930,G4931);
  nor NOR2_1549(G4989,G1301,G4932);
  nor NOR2_1550(G4993,G4935,G4870);
  nor NOR2_1551(G4997,G4938,G4875);
  nor NOR2_1552(G5001,G4941,G4880);
  nor NOR2_1553(G5005,G4944,G4885);
  nor NOR2_1554(G5009,G4893,G4947);
  nor NOR2_1555(G5010,G4947,G4890);
  nor NOR2_1556(G5011,G4951,G4952);
  nor NOR2_1557(G5014,G4953,G866);
  nor NOR2_1558(G5018,G4902,G4956);
  nor NOR2_1559(G5019,G4956,G914);
  nor NOR2_1560(G5020,G4776,G4956);
  nor NOR2_1561(G5023,G4960,G4961);
  nor NOR2_1562(G5026,G4965,G4962);
  nor NOR2_1563(G5030,G4914,G4968);
  nor NOR2_1564(G5031,G4968,G4911);
  nor NOR2_1565(G5032,G4972,G4973);
  nor NOR2_1566(G5035,G4974,G1109);
  nor NOR2_1567(G5039,G4923,G4977);
  nor NOR2_1568(G5040,G4977,G1157);
  nor NOR2_1569(G5041,G4797,G4977);
  nor NOR2_1570(G5044,G4981,G4982);
  nor NOR2_1571(G5047,G4986,G4983);
  nor NOR2_1572(G5051,G1301,G4989);
  nor NOR2_1573(G5052,G4989,G4932);
  nor NOR2_1574(G5053,G4935,G4993);
  nor NOR2_1575(G5054,G4993,G4870);
  nor NOR2_1576(G5055,G4938,G4997);
  nor NOR2_1577(G5056,G4997,G4875);
  nor NOR2_1578(G5057,G4941,G5001);
  nor NOR2_1579(G5058,G5001,G4880);
  nor NOR2_1580(G5059,G4944,G5005);
  nor NOR2_1581(G5060,G5005,G4885);
  nor NOR2_1582(G5061,G5009,G5010);
  nor NOR2_1583(G5064,G5011,G818);
  nor NOR2_1584(G5068,G4953,G5014);
  nor NOR2_1585(G5069,G5014,G866);
  nor NOR2_1586(G5070,G4834,G5014);
  nor NOR2_1587(G5073,G5018,G5019);
  nor NOR2_1588(G5076,G5023,G5020);
  nor NOR2_1589(G5080,G4965,G5026);
  nor NOR2_1590(G5081,G5026,G4962);
  nor NOR2_1591(G5082,G5030,G5031);
  nor NOR2_1592(G5085,G5032,G1061);
  nor NOR2_1593(G5089,G4974,G5035);
  nor NOR2_1594(G5090,G5035,G1109);
  nor NOR2_1595(G5091,G4855,G5035);
  nor NOR2_1596(G5094,G5039,G5040);
  nor NOR2_1597(G5097,G5044,G5041);
  nor NOR2_1598(G5101,G4986,G5047);
  nor NOR2_1599(G5102,G5047,G4983);
  nor NOR2_1600(G5103,G5051,G5052);
  nor NOR2_1601(G5106,G5053,G5054);
  nor NOR2_1602(G5109,G5055,G5056);
  nor NOR2_1603(G5112,G5057,G5058);
  nor NOR2_1604(G5115,G5059,G5060);
  nor NOR2_1605(G5118,G5061,G770);
  nor NOR2_1606(G5122,G5011,G5064);
  nor NOR2_1607(G5123,G5064,G818);
  nor NOR2_1608(G5124,G4896,G5064);
  nor NOR2_1609(G5127,G5068,G5069);
  nor NOR2_1610(G5130,G5073,G5070);
  nor NOR2_1611(G5134,G5023,G5076);
  nor NOR2_1612(G5135,G5076,G5020);
  nor NOR2_1613(G5136,G5080,G5081);
  nor NOR2_1614(G5139,G5082,G1013);
  nor NOR2_1615(G5143,G5032,G5085);
  nor NOR2_1616(G5144,G5085,G1061);
  nor NOR2_1617(G5145,G4917,G5085);
  nor NOR2_1618(G5148,G5089,G5090);
  nor NOR2_1619(G5151,G5094,G5091);
  nor NOR2_1620(G5155,G5044,G5097);
  nor NOR2_1621(G5156,G5097,G5041);
  nor NOR2_1622(G5157,G5101,G5102);
  nor NOR2_1623(G5160,G5103,G1256);
  nor NOR2_1624(G5164,G5106,G578);
  nor NOR2_1625(G5168,G5109,G626);
  nor NOR2_1626(G5172,G5112,G674);
  nor NOR2_1627(G5176,G5115,G722);
  nor NOR2_1628(G5180,G5061,G5118);
  nor NOR2_1629(G5181,G5118,G770);
  nor NOR2_1630(G5182,G4947,G5118);
  nor NOR2_1631(G5185,G5122,G5123);
  nor NOR2_1632(G5188,G5127,G5124);
  nor NOR2_1633(G5192,G5073,G5130);
  nor NOR2_1634(G5193,G5130,G5070);
  nor NOR2_1635(G5194,G5134,G5135);
  nor NOR2_1636(G5197,G5136,G965);
  nor NOR2_1637(G5201,G5082,G5139);
  nor NOR2_1638(G5202,G5139,G1013);
  nor NOR2_1639(G5203,G4968,G5139);
  nor NOR2_1640(G5206,G5143,G5144);
  nor NOR2_1641(G5209,G5148,G5145);
  nor NOR2_1642(G5213,G5094,G5151);
  nor NOR2_1643(G5214,G5151,G5091);
  nor NOR2_1644(G5215,G5155,G5156);
  nor NOR2_1645(G5218,G5157,G1208);
  nor NOR2_1646(G5222,G5103,G5160);
  nor NOR2_1647(G5223,G5160,G1256);
  nor NOR2_1648(G5224,G4989,G5160);
  nor NOR2_1649(G5227,G5106,G5164);
  nor NOR2_1650(G5228,G5164,G578);
  nor NOR2_1651(G5229,G4993,G5164);
  nor NOR2_1652(G5232,G5109,G5168);
  nor NOR2_1653(G5233,G5168,G626);
  nor NOR2_1654(G5234,G4997,G5168);
  nor NOR2_1655(G5237,G5112,G5172);
  nor NOR2_1656(G5238,G5172,G674);
  nor NOR2_1657(G5239,G5001,G5172);
  nor NOR2_1658(G5242,G5115,G5176);
  nor NOR2_1659(G5243,G5176,G722);
  nor NOR2_1660(G5244,G5005,G5176);
  nor NOR2_1661(G5247,G5180,G5181);
  nor NOR2_1662(G5250,G5185,G5182);
  nor NOR2_1663(G5254,G5127,G5188);
  nor NOR2_1664(G5255,G5188,G5124);
  nor NOR2_1665(G5256,G5192,G5193);
  nor NOR2_1666(G5259,G5194,G917);
  nor NOR2_1667(G5263,G5136,G5197);
  nor NOR2_1668(G5264,G5197,G965);
  nor NOR2_1669(G5265,G5026,G5197);
  nor NOR2_1670(G5268,G5201,G5202);
  nor NOR2_1671(G5271,G5206,G5203);
  nor NOR2_1672(G5275,G5148,G5209);
  nor NOR2_1673(G5276,G5209,G5145);
  nor NOR2_1674(G5277,G5213,G5214);
  nor NOR2_1675(G5280,G5215,G1160);
  nor NOR2_1676(G5284,G5157,G5218);
  nor NOR2_1677(G5285,G5218,G1208);
  nor NOR2_1678(G5286,G5047,G5218);
  nor NOR2_1679(G5289,G5222,G5223);
  nor NOR2_1680(G5292,G1304,G5224);
  nor NOR2_1681(G5296,G5232,G5233);
  nor NOR2_1682(G5299,G5237,G5238);
  nor NOR2_1683(G5302,G5242,G5243);
  nor NOR2_1684(G5305,G5247,G5244);
  nor NOR2_1685(G5309,G5185,G5250);
  nor NOR2_1686(G5310,G5250,G5182);
  nor NOR2_1687(G5311,G5254,G5255);
  nor NOR2_1688(G5314,G5256,G869);
  nor NOR2_1689(G5318,G5194,G5259);
  nor NOR2_1690(G5319,G5259,G917);
  nor NOR2_1691(G5320,G5076,G5259);
  nor NOR2_1692(G5323,G5263,G5264);
  nor NOR2_1693(G5326,G5268,G5265);
  nor NOR2_1694(G5330,G5206,G5271);
  nor NOR2_1695(G5331,G5271,G5203);
  nor NOR2_1696(G5332,G5275,G5276);
  nor NOR2_1697(G5335,G5277,G1112);
  nor NOR2_1698(G5339,G5215,G5280);
  nor NOR2_1699(G5340,G5280,G1160);
  nor NOR2_1700(G5341,G5097,G5280);
  nor NOR2_1701(G5344,G5284,G5285);
  nor NOR2_1702(G5347,G5289,G5286);
  nor NOR2_1703(G5351,G1304,G5292);
  nor NOR2_1704(G5352,G5292,G5224);
  nor NOR2_1705(G5353,G5296,G5229);
  nor NOR2_1706(G5357,G5299,G5234);
  nor NOR2_1707(G5361,G5302,G5239);
  nor NOR2_1708(G5365,G5247,G5305);
  nor NOR2_1709(G5366,G5305,G5244);
  nor NOR2_1710(G5367,G5309,G5310);
  nor NOR2_1711(G5370,G5311,G821);
  nor NOR2_1712(G5374,G5256,G5314);
  nor NOR2_1713(G5375,G5314,G869);
  nor NOR2_1714(G5376,G5130,G5314);
  nor NOR2_1715(G5379,G5318,G5319);
  nor NOR2_1716(G5382,G5323,G5320);
  nor NOR2_1717(G5386,G5268,G5326);
  nor NOR2_1718(G5387,G5326,G5265);
  nor NOR2_1719(G5388,G5330,G5331);
  nor NOR2_1720(G5391,G5332,G1064);
  nor NOR2_1721(G5395,G5277,G5335);
  nor NOR2_1722(G5396,G5335,G1112);
  nor NOR2_1723(G5397,G5151,G5335);
  nor NOR2_1724(G5400,G5339,G5340);
  nor NOR2_1725(G5403,G5344,G5341);
  nor NOR2_1726(G5407,G5289,G5347);
  nor NOR2_1727(G5408,G5347,G5286);
  nor NOR2_1728(G5409,G5351,G5352);
  nor NOR2_1729(G5412,G5296,G5353);
  nor NOR2_1730(G5413,G5353,G5229);
  nor NOR2_1731(G5414,G5299,G5357);
  nor NOR2_1732(G5415,G5357,G5234);
  nor NOR2_1733(G5416,G5302,G5361);
  nor NOR2_1734(G5417,G5361,G5239);
  nor NOR2_1735(G5418,G5365,G5366);
  nor NOR2_1736(G5421,G5367,G773);
  nor NOR2_1737(G5425,G5311,G5370);
  nor NOR2_1738(G5426,G5370,G821);
  nor NOR2_1739(G5427,G5188,G5370);
  nor NOR2_1740(G5430,G5374,G5375);
  nor NOR2_1741(G5433,G5379,G5376);
  nor NOR2_1742(G5437,G5323,G5382);
  nor NOR2_1743(G5438,G5382,G5320);
  nor NOR2_1744(G5439,G5386,G5387);
  nor NOR2_1745(G5442,G5388,G1016);
  nor NOR2_1746(G5446,G5332,G5391);
  nor NOR2_1747(G5447,G5391,G1064);
  nor NOR2_1748(G5448,G5209,G5391);
  nor NOR2_1749(G5451,G5395,G5396);
  nor NOR2_1750(G5454,G5400,G5397);
  nor NOR2_1751(G5458,G5344,G5403);
  nor NOR2_1752(G5459,G5403,G5341);
  nor NOR2_1753(G5460,G5407,G5408);
  nor NOR2_1754(G5463,G5409,G1259);
  nor NOR2_1755(G5467,G5412,G5413);
  nor NOR2_1756(G5470,G5414,G5415);
  nor NOR2_1757(G5473,G5416,G5417);
  nor NOR2_1758(G5476,G5418,G725);
  nor NOR2_1759(G5480,G5367,G5421);
  nor NOR2_1760(G5481,G5421,G773);
  nor NOR2_1761(G5482,G5250,G5421);
  nor NOR2_1762(G5485,G5425,G5426);
  nor NOR2_1763(G5488,G5430,G5427);
  nor NOR2_1764(G5492,G5379,G5433);
  nor NOR2_1765(G5493,G5433,G5376);
  nor NOR2_1766(G5494,G5437,G5438);
  nor NOR2_1767(G5497,G5439,G968);
  nor NOR2_1768(G5501,G5388,G5442);
  nor NOR2_1769(G5502,G5442,G1016);
  nor NOR2_1770(G5503,G5271,G5442);
  nor NOR2_1771(G5506,G5446,G5447);
  nor NOR2_1772(G5509,G5451,G5448);
  nor NOR2_1773(G5513,G5400,G5454);
  nor NOR2_1774(G5514,G5454,G5397);
  nor NOR2_1775(G5515,G5458,G5459);
  nor NOR2_1776(G5518,G5460,G1211);
  nor NOR2_1777(G5522,G5409,G5463);
  nor NOR2_1778(G5523,G5463,G1259);
  nor NOR2_1779(G5524,G5292,G5463);
  nor NOR2_1780(G5527,G5467,G581);
  nor NOR2_1781(G5531,G5470,G629);
  nor NOR2_1782(G5535,G5473,G677);
  nor NOR2_1783(G5539,G5418,G5476);
  nor NOR2_1784(G5540,G5476,G725);
  nor NOR2_1785(G5541,G5305,G5476);
  nor NOR2_1786(G5544,G5480,G5481);
  nor NOR2_1787(G5547,G5485,G5482);
  nor NOR2_1788(G5551,G5430,G5488);
  nor NOR2_1789(G5552,G5488,G5427);
  nor NOR2_1790(G5553,G5492,G5493);
  nor NOR2_1791(G5556,G5494,G920);
  nor NOR2_1792(G5560,G5439,G5497);
  nor NOR2_1793(G5561,G5497,G968);
  nor NOR2_1794(G5562,G5326,G5497);
  nor NOR2_1795(G5565,G5501,G5502);
  nor NOR2_1796(G5568,G5506,G5503);
  nor NOR2_1797(G5572,G5451,G5509);
  nor NOR2_1798(G5573,G5509,G5448);
  nor NOR2_1799(G5574,G5513,G5514);
  nor NOR2_1800(G5577,G5515,G1163);
  nor NOR2_1801(G5581,G5460,G5518);
  nor NOR2_1802(G5582,G5518,G1211);
  nor NOR2_1803(G5583,G5347,G5518);
  nor NOR2_1804(G5586,G5522,G5523);
  nor NOR2_1805(G5589,G1307,G5524);
  nor NOR2_1806(G5593,G5467,G5527);
  nor NOR2_1807(G5594,G5527,G581);
  nor NOR2_1808(G5595,G5353,G5527);
  nor NOR2_1809(G5598,G5470,G5531);
  nor NOR2_1810(G5599,G5531,G629);
  nor NOR2_1811(G5600,G5357,G5531);
  nor NOR2_1812(G5603,G5473,G5535);
  nor NOR2_1813(G5604,G5535,G677);
  nor NOR2_1814(G5605,G5361,G5535);
  nor NOR2_1815(G5608,G5539,G5540);
  nor NOR2_1816(G5611,G5544,G5541);
  nor NOR2_1817(G5615,G5485,G5547);
  nor NOR2_1818(G5616,G5547,G5482);
  nor NOR2_1819(G5617,G5551,G5552);
  nor NOR2_1820(G5620,G5553,G872);
  nor NOR2_1821(G5624,G5494,G5556);
  nor NOR2_1822(G5625,G5556,G920);
  nor NOR2_1823(G5626,G5382,G5556);
  nor NOR2_1824(G5629,G5560,G5561);
  nor NOR2_1825(G5632,G5565,G5562);
  nor NOR2_1826(G5636,G5506,G5568);
  nor NOR2_1827(G5637,G5568,G5503);
  nor NOR2_1828(G5638,G5572,G5573);
  nor NOR2_1829(G5641,G5574,G1115);
  nor NOR2_1830(G5645,G5515,G5577);
  nor NOR2_1831(G5646,G5577,G1163);
  nor NOR2_1832(G5647,G5403,G5577);
  nor NOR2_1833(G5650,G5581,G5582);
  nor NOR2_1834(G5653,G5586,G5583);
  nor NOR2_1835(G5657,G1307,G5589);
  nor NOR2_1836(G5658,G5589,G5524);
  nor NOR2_1837(G5659,G5598,G5599);
  nor NOR2_1838(G5662,G5603,G5604);
  nor NOR2_1839(G5665,G5608,G5605);
  nor NOR2_1840(G5669,G5544,G5611);
  nor NOR2_1841(G5670,G5611,G5541);
  nor NOR2_1842(G5671,G5615,G5616);
  nor NOR2_1843(G5674,G5617,G824);
  nor NOR2_1844(G5678,G5553,G5620);
  nor NOR2_1845(G5679,G5620,G872);
  nor NOR2_1846(G5680,G5433,G5620);
  nor NOR2_1847(G5683,G5624,G5625);
  nor NOR2_1848(G5686,G5629,G5626);
  nor NOR2_1849(G5690,G5565,G5632);
  nor NOR2_1850(G5691,G5632,G5562);
  nor NOR2_1851(G5692,G5636,G5637);
  nor NOR2_1852(G5695,G5638,G1067);
  nor NOR2_1853(G5699,G5574,G5641);
  nor NOR2_1854(G5700,G5641,G1115);
  nor NOR2_1855(G5701,G5454,G5641);
  nor NOR2_1856(G5704,G5645,G5646);
  nor NOR2_1857(G5707,G5650,G5647);
  nor NOR2_1858(G5711,G5586,G5653);
  nor NOR2_1859(G5712,G5653,G5583);
  nor NOR2_1860(G5713,G5657,G5658);
  nor NOR2_1861(G5716,G5659,G5595);
  nor NOR2_1862(G5720,G5662,G5600);
  nor NOR2_1863(G5724,G5608,G5665);
  nor NOR2_1864(G5725,G5665,G5605);
  nor NOR2_1865(G5726,G5669,G5670);
  nor NOR2_1866(G5729,G5671,G776);
  nor NOR2_1867(G5733,G5617,G5674);
  nor NOR2_1868(G5734,G5674,G824);
  nor NOR2_1869(G5735,G5488,G5674);
  nor NOR2_1870(G5738,G5678,G5679);
  nor NOR2_1871(G5741,G5683,G5680);
  nor NOR2_1872(G5745,G5629,G5686);
  nor NOR2_1873(G5746,G5686,G5626);
  nor NOR2_1874(G5747,G5690,G5691);
  nor NOR2_1875(G5750,G5692,G1019);
  nor NOR2_1876(G5754,G5638,G5695);
  nor NOR2_1877(G5755,G5695,G1067);
  nor NOR2_1878(G5756,G5509,G5695);
  nor NOR2_1879(G5759,G5699,G5700);
  nor NOR2_1880(G5762,G5704,G5701);
  nor NOR2_1881(G5766,G5650,G5707);
  nor NOR2_1882(G5767,G5707,G5647);
  nor NOR2_1883(G5768,G5711,G5712);
  nor NOR2_1884(G5771,G5659,G5716);
  nor NOR2_1885(G5772,G5716,G5595);
  nor NOR2_1886(G5773,G5662,G5720);
  nor NOR2_1887(G5774,G5720,G5600);
  nor NOR2_1888(G5775,G5724,G5725);
  nor NOR2_1889(G5778,G5726,G728);
  nor NOR2_1890(G5782,G5671,G5729);
  nor NOR2_1891(G5783,G5729,G776);
  nor NOR2_1892(G5784,G5547,G5729);
  nor NOR2_1893(G5787,G5733,G5734);
  nor NOR2_1894(G5790,G5738,G5735);
  nor NOR2_1895(G5794,G5683,G5741);
  nor NOR2_1896(G5795,G5741,G5680);
  nor NOR2_1897(G5796,G5745,G5746);
  nor NOR2_1898(G5799,G5747,G971);
  nor NOR2_1899(G5803,G5692,G5750);
  nor NOR2_1900(G5804,G5750,G1019);
  nor NOR2_1901(G5805,G5568,G5750);
  nor NOR2_1902(G5808,G5754,G5755);
  nor NOR2_1903(G5811,G5759,G5756);
  nor NOR2_1904(G5815,G5704,G5762);
  nor NOR2_1905(G5816,G5762,G5701);
  nor NOR2_1906(G5817,G5766,G5767);
  nor NOR2_1907(G5820,G5771,G5772);
  nor NOR2_1908(G5823,G5773,G5774);
  nor NOR2_1909(G5826,G5775,G680);
  nor NOR2_1910(G5830,G5726,G5778);
  nor NOR2_1911(G5831,G5778,G728);
  nor NOR2_1912(G5832,G5611,G5778);
  nor NOR2_1913(G5835,G5782,G5783);
  nor NOR2_1914(G5838,G5787,G5784);
  nor NOR2_1915(G5842,G5738,G5790);
  nor NOR2_1916(G5843,G5790,G5735);
  nor NOR2_1917(G5844,G5794,G5795);
  nor NOR2_1918(G5847,G5796,G923);
  nor NOR2_1919(G5851,G5747,G5799);
  nor NOR2_1920(G5852,G5799,G971);
  nor NOR2_1921(G5853,G5632,G5799);
  nor NOR2_1922(G5856,G5803,G5804);
  nor NOR2_1923(G5859,G5808,G5805);
  nor NOR2_1924(G5863,G5759,G5811);
  nor NOR2_1925(G5864,G5811,G5756);
  nor NOR2_1926(G5865,G5815,G5816);
  nor NOR2_1927(G5868,G5820,G584);
  nor NOR2_1928(G5872,G5823,G632);
  nor NOR2_1929(G5876,G5775,G5826);
  nor NOR2_1930(G5877,G5826,G680);
  nor NOR2_1931(G5878,G5665,G5826);
  nor NOR2_1932(G5881,G5830,G5831);
  nor NOR2_1933(G5884,G5835,G5832);
  nor NOR2_1934(G5888,G5787,G5838);
  nor NOR2_1935(G5889,G5838,G5784);
  nor NOR2_1936(G5890,G5842,G5843);
  nor NOR2_1937(G5893,G5844,G875);
  nor NOR2_1938(G5897,G5796,G5847);
  nor NOR2_1939(G5898,G5847,G923);
  nor NOR2_1940(G5899,G5686,G5847);
  nor NOR2_1941(G5902,G5851,G5852);
  nor NOR2_1942(G5905,G5856,G5853);
  nor NOR2_1943(G5909,G5808,G5859);
  nor NOR2_1944(G5910,G5859,G5805);
  nor NOR2_1945(G5911,G5863,G5864);
  nor NOR2_1946(G5914,G5820,G5868);
  nor NOR2_1947(G5915,G5868,G584);
  nor NOR2_1948(G5916,G5716,G5868);
  nor NOR2_1949(G5919,G5823,G5872);
  nor NOR2_1950(G5920,G5872,G632);
  nor NOR2_1951(G5921,G5720,G5872);
  nor NOR2_1952(G5924,G5876,G5877);
  nor NOR2_1953(G5927,G5881,G5878);
  nor NOR2_1954(G5931,G5835,G5884);
  nor NOR2_1955(G5932,G5884,G5832);
  nor NOR2_1956(G5933,G5888,G5889);
  nor NOR2_1957(G5936,G5890,G827);
  nor NOR2_1958(G5940,G5844,G5893);
  nor NOR2_1959(G5941,G5893,G875);
  nor NOR2_1960(G5942,G5741,G5893);
  nor NOR2_1961(G5945,G5897,G5898);
  nor NOR2_1962(G5948,G5902,G5899);
  nor NOR2_1963(G5952,G5856,G5905);
  nor NOR2_1964(G5953,G5905,G5853);
  nor NOR2_1965(G5954,G5909,G5910);
  nor NOR2_1966(G5957,G5919,G5920);
  nor NOR2_1967(G5960,G5924,G5921);
  nor NOR2_1968(G5964,G5881,G5927);
  nor NOR2_1969(G5965,G5927,G5878);
  nor NOR2_1970(G5966,G5931,G5932);
  nor NOR2_1971(G5969,G5933,G779);
  nor NOR2_1972(G5973,G5890,G5936);
  nor NOR2_1973(G5974,G5936,G827);
  nor NOR2_1974(G5975,G5790,G5936);
  nor NOR2_1975(G5978,G5940,G5941);
  nor NOR2_1976(G5981,G5945,G5942);
  nor NOR2_1977(G5985,G5902,G5948);
  nor NOR2_1978(G5986,G5948,G5899);
  nor NOR2_1979(G5987,G5952,G5953);
  nor NOR2_1980(G5990,G5957,G5916);
  nor NOR2_1981(G5994,G5924,G5960);
  nor NOR2_1982(G5995,G5960,G5921);
  nor NOR2_1983(G5996,G5964,G5965);
  nor NOR2_1984(G5999,G5966,G731);
  nor NOR2_1985(G6003,G5933,G5969);
  nor NOR2_1986(G6004,G5969,G779);
  nor NOR2_1987(G6005,G5838,G5969);
  nor NOR2_1988(G6008,G5973,G5974);
  nor NOR2_1989(G6011,G5978,G5975);
  nor NOR2_1990(G6015,G5945,G5981);
  nor NOR2_1991(G6016,G5981,G5942);
  nor NOR2_1992(G6017,G5985,G5986);
  nor NOR2_1993(G6020,G5957,G5990);
  nor NOR2_1994(G6021,G5990,G5916);
  nor NOR2_1995(G6022,G5994,G5995);
  nor NOR2_1996(G6025,G5996,G683);
  nor NOR2_1997(G6029,G5966,G5999);
  nor NOR2_1998(G6030,G5999,G731);
  nor NOR2_1999(G6031,G5884,G5999);
  nor NOR2_2000(G6034,G6003,G6004);
  nor NOR2_2001(G6037,G6008,G6005);
  nor NOR2_2002(G6041,G5978,G6011);
  nor NOR2_2003(G6042,G6011,G5975);
  nor NOR2_2004(G6043,G6015,G6016);
  nor NOR2_2005(G6046,G6020,G6021);
  nor NOR2_2006(G6049,G6022,G635);
  nor NOR2_2007(G6053,G5996,G6025);
  nor NOR2_2008(G6054,G6025,G683);
  nor NOR2_2009(G6055,G5927,G6025);
  nor NOR2_2010(G6058,G6029,G6030);
  nor NOR2_2011(G6061,G6034,G6031);
  nor NOR2_2012(G6065,G6008,G6037);
  nor NOR2_2013(G6066,G6037,G6005);
  nor NOR2_2014(G6067,G6041,G6042);
  nor NOR2_2015(G6070,G6046,G587);
  nor NOR2_2016(G6074,G6022,G6049);
  nor NOR2_2017(G6075,G6049,G635);
  nor NOR2_2018(G6076,G5960,G6049);
  nor NOR2_2019(G6079,G6053,G6054);
  nor NOR2_2020(G6082,G6058,G6055);
  nor NOR2_2021(G6086,G6034,G6061);
  nor NOR2_2022(G6087,G6061,G6031);
  nor NOR2_2023(G6088,G6065,G6066);
  nor NOR2_2024(G6091,G6046,G6070);
  nor NOR2_2025(G6092,G6070,G587);
  nor NOR2_2026(G6093,G5990,G6070);
  nor NOR2_2027(G6096,G6074,G6075);
  nor NOR2_2028(G6099,G6079,G6076);
  nor NOR2_2029(G6103,G6058,G6082);
  nor NOR2_2030(G6104,G6082,G6055);
  nor NOR2_2031(G6105,G6086,G6087);
  nor NOR2_2032(G6108,G6096,G6093);
  nor NOR2_2033(G6112,G6079,G6099);
  nor NOR2_2034(G6113,G6099,G6076);
  nor NOR2_2035(G6114,G6103,G6104);
  nor NOR2_2036(G6117,G6096,G6108);
  nor NOR2_2037(G6118,G6108,G6093);
  nor NOR2_2038(G6119,G6112,G6113);
  nor NOR2_2039(G6122,G6117,G6118);
  not NOT_30(G6125,G6122);
  nor NOR2_2040(G6129,G6122,G6125);
  not NOT_31(G6130,G6125);
  nor NOR2_2041(G6131,G6108,G6125);
  nor NOR2_2042(G6134,G6119,G6131);
  nor NOR2_2043(G6138,G6119,G6134);
  nor NOR2_2044(G6139,G6134,G6131);
  nor NOR2_2045(G6140,G6099,G6134);
  nor NOR2_2046(G6143,G6114,G6140);
  nor NOR2_2047(G6147,G6114,G6143);
  nor NOR2_2048(G6148,G6143,G6140);
  nor NOR2_2049(G6149,G6082,G6143);
  nor NOR2_2050(G6152,G6105,G6149);
  nor NOR2_2051(G6156,G6105,G6152);
  nor NOR2_2052(G6157,G6152,G6149);
  nor NOR2_2053(G6158,G6061,G6152);
  nor NOR2_2054(G6161,G6088,G6158);
  nor NOR2_2055(G6165,G6088,G6161);
  nor NOR2_2056(G6166,G6161,G6158);
  nor NOR2_2057(G6167,G6037,G6161);
  nor NOR2_2058(G6170,G6067,G6167);
  nor NOR2_2059(G6174,G6067,G6170);
  nor NOR2_2060(G6175,G6170,G6167);
  nor NOR2_2061(G6176,G6011,G6170);
  nor NOR2_2062(G6179,G6043,G6176);
  nor NOR2_2063(G6183,G6043,G6179);
  nor NOR2_2064(G6184,G6179,G6176);
  nor NOR2_2065(G6185,G5981,G6179);
  nor NOR2_2066(G6188,G6017,G6185);
  nor NOR2_2067(G6192,G6017,G6188);
  nor NOR2_2068(G6193,G6188,G6185);
  nor NOR2_2069(G6194,G5948,G6188);
  nor NOR2_2070(G6197,G5987,G6194);
  nor NOR2_2071(G6201,G5987,G6197);
  nor NOR2_2072(G6202,G6197,G6194);
  nor NOR2_2073(G6203,G5905,G6197);
  nor NOR2_2074(G6206,G5954,G6203);
  nor NOR2_2075(G6210,G5954,G6206);
  nor NOR2_2076(G6211,G6206,G6203);
  nor NOR2_2077(G6212,G5859,G6206);
  nor NOR2_2078(G6215,G5911,G6212);
  nor NOR2_2079(G6219,G5911,G6215);
  nor NOR2_2080(G6220,G6215,G6212);
  nor NOR2_2081(G6221,G5811,G6215);
  nor NOR2_2082(G6224,G5865,G6221);
  nor NOR2_2083(G6228,G5865,G6224);
  nor NOR2_2084(G6229,G6224,G6221);
  nor NOR2_2085(G6230,G5762,G6224);
  nor NOR2_2086(G6233,G5817,G6230);
  nor NOR2_2087(G6237,G5817,G6233);
  nor NOR2_2088(G6238,G6233,G6230);
  nor NOR2_2089(G6239,G5707,G6233);
  nor NOR2_2090(G6242,G5768,G6239);
  nor NOR2_2091(G6246,G5768,G6242);
  nor NOR2_2092(G6247,G6242,G6239);
  nor NOR2_2093(G6248,G5653,G6242);
  nor NOR2_2094(G6251,G5713,G6248);
  nor NOR2_2095(G6255,G5713,G6251);
  nor NOR2_2096(G6256,G6251,G6248);
  and AND2_255(G6257,G1,G17);
  nor NOR2_2097(G6258,G1505,G1506);
  nor NOR2_2098(G6259,G1822,G1823);
  nor NOR2_2099(G6260,G2146,G2147);
  nor NOR2_2100(G6261,G2472,G2473);
  nor NOR2_2101(G6262,G2801,G2802);
  nor NOR2_2102(G6263,G3134,G3135);
  nor NOR2_2103(G6264,G3472,G3473);
  nor NOR2_2104(G6265,G3817,G3818);
  nor NOR2_2105(G6266,G4164,G4165);
  nor NOR2_2106(G6267,G4514,G4515);
  nor NOR2_2107(G6268,G4868,G4869);
  nor NOR2_2108(G6269,G5227,G5228);
  nor NOR2_2109(G6270,G5593,G5594);
  nor NOR2_2110(G6271,G5914,G5915);
  nor NOR2_2111(G6272,G6091,G6092);
  nor NOR2_2112(G6273,G6129,G6130);
  nor NOR2_2113(G6274,G6138,G6139);
  nor NOR2_2114(G6275,G6147,G6148);
  nor NOR2_2115(G6276,G6156,G6157);
  nor NOR2_2116(G6277,G6165,G6166);
  nor NOR2_2117(G6278,G6174,G6175);
  nor NOR2_2118(G6279,G6183,G6184);
  nor NOR2_2119(G6280,G6192,G6193);
  nor NOR2_2120(G6281,G6201,G6202);
  nor NOR2_2121(G6282,G6210,G6211);
  nor NOR2_2122(G6283,G6219,G6220);
  nor NOR2_2123(G6284,G6228,G6229);
  nor NOR2_2124(G6285,G6237,G6238);
  nor NOR2_2125(G6286,G6246,G6247);
  nor NOR2_2126(G6287,G5589,G6251);
  nor NOR2_2127(G6288,G6255,G6256);

endmodule
