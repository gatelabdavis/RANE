module c499(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,
  G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,
  G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,G481,G482,
  G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,
  G498,G499,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,G481,
  G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,
  G497,G498,G499;

  wire G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,
    G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,
    G175,G176,G177,G178,G179,G180,G181,G182,G183,G184,G185,G186,G189,G192,G195,
    G198,G201,G204,G207,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
    G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G247,
    G260,G273,G286,G299,G312,G325,G338,G339,G340,G341,G342,G343,G344,G345,G346,
    G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,G361,
    G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,
    G377,G378,G379,G380,G381,G382,G383,G384,G385,G386,G391,G396,G401,G406,G411,
    G416,G421,G426,G431,G436,G437,G438,G439,G440,G441,G442,G443,G444,G445,G446,
    G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,G461,
    G462,G463,G464,G465,G466,G467;

  xor XOR2_0(G146,G1,G2);
  xor XOR2_1(G147,G3,G4);
  xor XOR2_2(G148,G5,G6);
  xor XOR2_3(G149,G7,G8);
  xor XOR2_4(G150,G9,G10);
  xor XOR2_5(G151,G11,G12);
  xor XOR2_6(G152,G13,G14);
  xor XOR2_7(G153,G15,G16);
  xor XOR2_8(G154,G17,G18);
  xor XOR2_9(G155,G19,G20);
  xor XOR2_10(G156,G21,G22);
  xor XOR2_11(G157,G23,G24);
  xor XOR2_12(G158,G25,G26);
  xor XOR2_13(G159,G27,G28);
  xor XOR2_14(G160,G29,G30);
  xor XOR2_15(G161,G31,G32);
  and AND2_0(G162,G33,G41);
  and AND2_1(G163,G34,G41);
  and AND2_2(G164,G35,G41);
  and AND2_3(G165,G36,G41);
  and AND2_4(G166,G37,G41);
  and AND2_5(G167,G38,G41);
  and AND2_6(G168,G39,G41);
  and AND2_7(G169,G40,G41);
  xor XOR2_16(G170,G1,G5);
  xor XOR2_17(G171,G9,G13);
  xor XOR2_18(G172,G2,G6);
  xor XOR2_19(G173,G10,G14);
  xor XOR2_20(G174,G3,G7);
  xor XOR2_21(G175,G11,G15);
  xor XOR2_22(G176,G4,G8);
  xor XOR2_23(G177,G12,G16);
  xor XOR2_24(G178,G17,G21);
  xor XOR2_25(G179,G25,G29);
  xor XOR2_26(G180,G18,G22);
  xor XOR2_27(G181,G26,G30);
  xor XOR2_28(G182,G19,G23);
  xor XOR2_29(G183,G27,G31);
  xor XOR2_30(G184,G20,G24);
  xor XOR2_31(G185,G28,G32);
  xor XOR2_32(G186,G146,G147);
  xor XOR2_33(G189,G148,G149);
  xor XOR2_34(G192,G150,G151);
  xor XOR2_35(G195,G152,G153);
  xor XOR2_36(G198,G154,G155);
  xor XOR2_37(G201,G156,G157);
  xor XOR2_38(G204,G158,G159);
  xor XOR2_39(G207,G160,G161);
  xor XOR2_40(G210,G170,G171);
  xor XOR2_41(G211,G172,G173);
  xor XOR2_42(G212,G174,G175);
  xor XOR2_43(G213,G176,G177);
  xor XOR2_44(G214,G178,G179);
  xor XOR2_45(G215,G180,G181);
  xor XOR2_46(G216,G182,G183);
  xor XOR2_47(G217,G184,G185);
  xor XOR2_48(G218,G186,G189);
  xor XOR2_49(G219,G192,G195);
  xor XOR2_50(G220,G186,G192);
  xor XOR2_51(G221,G189,G195);
  xor XOR2_52(G222,G198,G201);
  xor XOR2_53(G223,G204,G207);
  xor XOR2_54(G224,G198,G204);
  xor XOR2_55(G225,G201,G207);
  xor XOR2_56(G226,G162,G222);
  xor XOR2_57(G227,G163,G223);
  xor XOR2_58(G228,G164,G224);
  xor XOR2_59(G229,G165,G225);
  xor XOR2_60(G230,G166,G218);
  xor XOR2_61(G231,G167,G219);
  xor XOR2_62(G232,G168,G220);
  xor XOR2_63(G233,G169,G221);
  xor XOR2_64(G234,G210,G226);
  xor XOR2_65(G247,G211,G227);
  xor XOR2_66(G260,G212,G228);
  xor XOR2_67(G273,G213,G229);
  xor XOR2_68(G286,G214,G230);
  xor XOR2_69(G299,G215,G231);
  xor XOR2_70(G312,G216,G232);
  xor XOR2_71(G325,G217,G233);
  not NOT_0(G338,G234);
  not NOT_1(G339,G247);
  not NOT_2(G340,G260);
  not NOT_3(G341,G234);
  not NOT_4(G342,G247);
  not NOT_5(G343,G273);
  not NOT_6(G344,G234);
  not NOT_7(G345,G260);
  not NOT_8(G346,G273);
  not NOT_9(G347,G247);
  not NOT_10(G348,G260);
  not NOT_11(G349,G273);
  not NOT_12(G350,G299);
  not NOT_13(G351,G325);
  not NOT_14(G352,G299);
  not NOT_15(G353,G312);
  not NOT_16(G354,G286);
  not NOT_17(G355,G325);
  not NOT_18(G356,G286);
  not NOT_19(G357,G312);
  not NOT_20(G358,G286);
  not NOT_21(G359,G299);
  not NOT_22(G360,G312);
  not NOT_23(G361,G286);
  not NOT_24(G362,G299);
  not NOT_25(G363,G325);
  not NOT_26(G364,G286);
  not NOT_27(G365,G312);
  not NOT_28(G366,G325);
  not NOT_29(G367,G299);
  not NOT_30(G368,G312);
  not NOT_31(G369,G325);
  not NOT_32(G370,G247);
  not NOT_33(G371,G273);
  not NOT_34(G372,G247);
  not NOT_35(G373,G260);
  not NOT_36(G374,G234);
  not NOT_37(G375,G273);
  not NOT_38(G376,G234);
  not NOT_39(G377,G260);
  and AND4_0(G378,G338,G339,G340,G273);
  and AND4_1(G379,G341,G342,G260,G343);
  and AND4_2(G380,G344,G247,G345,G346);
  and AND4_3(G381,G234,G347,G348,G349);
  and AND4_4(G382,G358,G359,G360,G325);
  and AND4_5(G383,G361,G362,G312,G363);
  and AND4_6(G384,G364,G299,G365,G366);
  and AND4_7(G385,G286,G367,G368,G369);
  or OR4_0(G386,G378,G379,G380,G381);
  or OR4_1(G391,G382,G383,G384,G385);
  and AND5_0(G396,G286,G350,G312,G351,G386);
  and AND5_1(G401,G286,G352,G353,G325,G386);
  and AND5_2(G406,G354,G299,G312,G355,G386);
  and AND5_3(G411,G356,G299,G357,G325,G386);
  and AND5_4(G416,G234,G370,G260,G371,G391);
  and AND5_5(G421,G234,G372,G373,G273,G391);
  and AND5_6(G426,G374,G247,G260,G375,G391);
  and AND5_7(G431,G376,G247,G377,G273,G391);
  and AND2_8(G436,G234,G396);
  and AND2_9(G437,G247,G396);
  and AND2_10(G438,G260,G396);
  and AND2_11(G439,G273,G396);
  and AND2_12(G440,G234,G401);
  and AND2_13(G441,G247,G401);
  and AND2_14(G442,G260,G401);
  and AND2_15(G443,G273,G401);
  and AND2_16(G444,G234,G406);
  and AND2_17(G445,G247,G406);
  and AND2_18(G446,G260,G406);
  and AND2_19(G447,G273,G406);
  and AND2_20(G448,G234,G411);
  and AND2_21(G449,G247,G411);
  and AND2_22(G450,G260,G411);
  and AND2_23(G451,G273,G411);
  and AND2_24(G452,G286,G416);
  and AND2_25(G453,G299,G416);
  and AND2_26(G454,G312,G416);
  and AND2_27(G455,G325,G416);
  and AND2_28(G456,G286,G421);
  and AND2_29(G457,G299,G421);
  and AND2_30(G458,G312,G421);
  and AND2_31(G459,G325,G421);
  and AND2_32(G460,G286,G426);
  and AND2_33(G461,G299,G426);
  and AND2_34(G462,G312,G426);
  and AND2_35(G463,G325,G426);
  and AND2_36(G464,G286,G431);
  and AND2_37(G465,G299,G431);
  and AND2_38(G466,G312,G431);
  and AND2_39(G467,G325,G431);
  xor XOR2_72(G468,G1,G436);
  xor XOR2_73(G469,G2,G437);
  xor XOR2_74(G470,G3,G438);
  xor XOR2_75(G471,G4,G439);
  xor XOR2_76(G472,G5,G440);
  xor XOR2_77(G473,G6,G441);
  xor XOR2_78(G474,G7,G442);
  xor XOR2_79(G475,G8,G443);
  xor XOR2_80(G476,G9,G444);
  xor XOR2_81(G477,G10,G445);
  xor XOR2_82(G478,G11,G446);
  xor XOR2_83(G479,G12,G447);
  xor XOR2_84(G480,G13,G448);
  xor XOR2_85(G481,G14,G449);
  xor XOR2_86(G482,G15,G450);
  xor XOR2_87(G483,G16,G451);
  xor XOR2_88(G484,G17,G452);
  xor XOR2_89(G485,G18,G453);
  xor XOR2_90(G486,G19,G454);
  xor XOR2_91(G487,G20,G455);
  xor XOR2_92(G488,G21,G456);
  xor XOR2_93(G489,G22,G457);
  xor XOR2_94(G490,G23,G458);
  xor XOR2_95(G491,G24,G459);
  xor XOR2_96(G492,G25,G460);
  xor XOR2_97(G493,G26,G461);
  xor XOR2_98(G494,G27,G462);
  xor XOR2_99(G495,G28,G463);
  xor XOR2_100(G496,G29,G464);
  xor XOR2_101(G497,G30,G465);
  xor XOR2_102(G498,G31,G466);
  xor XOR2_103(G499,G32,G467);

endmodule
