// key=010110111

module s27_obf(CK, G0, G1, G2, G3, G17, keyinput);
input CK;
input G0;
input G1;
input G2;
input G3;
input [8:0] keyinput;
output G17;
wire G5;
wire G6;
wire G7;
wire G14;
wire G14_obf;
wire G13;
wire G13_obf;
wire G11;
wire G11_obf;
wire G15;
wire G15_obf;
wire G8;
wire G8_obf;
wire G16;
wire G16_obf;
wire G10;
wire G10_obf;
wire G12;
wire G12_obf;
wire G9;
wire G9_obf;
dff DFF_0(CK, G5, G10);
dff DFF_1(CK, G6, G11);
dff DFF_2(CK, G7, G13);
not NOT_1(G17, G11);
xnor tag0(G14, keyinput[0], G14_obf);
not NOT_0(G14_obf, G0);
xnor tag1(G13, keyinput[1], G13_obf);
nor NOR2_3(G13_obf, G2, G12);
xnor tag2(G11, keyinput[2], G11_obf);
nor NOR2_1(G11_obf, G5, G9);
xor tag3(G15, keyinput[3], G15_obf);
or OR2_0(G15_obf, G12, G8);
xnor tag4(G8, keyinput[4], G8_obf);
and AND2_0(G8_obf, G14, G6);
xnor tag5(G16, keyinput[5], G16_obf);
or OR2_1(G16_obf, G3, G8);
xor tag6(G10, keyinput[6], G10_obf);
nor NOR2_0(G10_obf, G14, G11);
xnor tag7(G12, keyinput[7], G12_obf);
nor NOR2_2(G12_obf, G1, G7);
xor tag8(G9, keyinput[8], G9_obf);
nand NAND2_0(G9_obf, G16, G15);
endmodule